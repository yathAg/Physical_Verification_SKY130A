* Example SPICE netlist netA.spice
*
.subckt cell4 A B C
.ends

.subckt cell2 A B C
.ends

.subckt cell3 A B C
.ends

.subckt test A B C
X1 A B C cell4
X2 A B A cell2
X3 C C A cell3
.ends
.end
