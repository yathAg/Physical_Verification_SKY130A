magic
tech sky130A
magscale 1 2
timestamp 1665771558
<< error_p >>
rect -29 222 29 228
rect -29 188 -17 222
rect -29 182 29 188
rect -125 -188 -67 -182
rect 67 -188 125 -182
rect -125 -222 -113 -188
rect 67 -222 79 -188
rect -125 -228 -67 -222
rect 67 -228 125 -222
<< pwell >>
rect -311 -360 311 360
<< nmos >>
rect -114 -150 -78 150
rect -18 -150 18 150
rect 78 -150 114 150
<< ndiff >>
rect -173 138 -114 150
rect -173 -138 -161 138
rect -127 -138 -114 138
rect -173 -150 -114 -138
rect -78 138 -18 150
rect -78 -138 -65 138
rect -31 -138 -18 138
rect -78 -150 -18 -138
rect 18 138 78 150
rect 18 -138 31 138
rect 65 -138 78 138
rect 18 -150 78 -138
rect 114 138 173 150
rect 114 -138 127 138
rect 161 -138 173 138
rect 114 -150 173 -138
<< ndiffc >>
rect -161 -138 -127 138
rect -65 -138 -31 138
rect 31 -138 65 138
rect 127 -138 161 138
<< psubdiff >>
rect -275 290 -179 324
rect 179 290 275 324
rect -275 228 -241 290
rect 241 228 275 290
rect -275 -290 -241 -228
rect 241 -290 275 -228
rect -275 -324 -179 -290
rect 179 -324 275 -290
<< psubdiffcont >>
rect -179 290 179 324
rect -275 -228 -241 228
rect 241 -228 275 228
rect -179 -324 179 -290
<< poly >>
rect -33 222 33 238
rect -33 188 -17 222
rect 17 188 33 222
rect -114 150 -78 176
rect -33 172 33 188
rect -18 150 18 172
rect 78 150 114 176
rect -114 -172 -78 -150
rect -129 -188 -63 -172
rect -18 -176 18 -150
rect 78 -172 114 -150
rect -129 -222 -113 -188
rect -79 -222 -63 -188
rect -129 -238 -63 -222
rect 63 -188 129 -172
rect 63 -222 79 -188
rect 113 -222 129 -188
rect 63 -238 129 -222
<< polycont >>
rect -17 188 17 222
rect -113 -222 -79 -188
rect 79 -222 113 -188
<< locali >>
rect -275 290 -179 324
rect 179 290 275 324
rect -275 228 -241 290
rect 241 228 275 290
rect -33 188 -17 222
rect 17 188 33 222
rect -161 138 -127 154
rect -161 -154 -127 -138
rect -65 138 -31 154
rect -65 -154 -31 -138
rect 31 138 65 154
rect 31 -154 65 -138
rect 127 138 161 154
rect 127 -154 161 -138
rect -129 -222 -113 -188
rect -79 -222 -63 -188
rect 63 -222 79 -188
rect 113 -222 129 -188
rect -275 -324 -241 -228
rect 241 -324 275 -228
<< viali >>
rect -17 188 17 222
rect -161 11 -127 121
rect -65 -121 -31 -11
rect 31 11 65 121
rect 127 -121 161 -11
rect -113 -222 -79 -188
rect 79 -222 113 -188
rect -241 -324 -179 -290
rect -179 -324 179 -290
rect 179 -324 241 -290
<< metal1 >>
rect -29 222 29 228
rect -29 188 -17 222
rect 17 188 29 222
rect -29 182 29 188
rect -167 121 -121 133
rect -167 11 -161 121
rect -127 11 -121 121
rect -167 -1 -121 11
rect 25 121 71 133
rect 25 11 31 121
rect 65 11 71 121
rect -71 -11 -25 1
rect 25 -1 71 11
rect -71 -121 -65 -11
rect -31 -121 -25 -11
rect -71 -133 -25 -121
rect 121 -11 167 1
rect 121 -121 127 -11
rect 161 -121 167 -11
rect 121 -133 167 -121
rect -125 -188 -67 -182
rect -125 -222 -113 -188
rect -79 -222 -67 -188
rect -125 -228 -67 -222
rect 67 -188 125 -182
rect 67 -222 79 -188
rect 113 -222 125 -188
rect 67 -228 125 -222
rect -253 -290 253 -284
rect -253 -324 -241 -290
rect 241 -324 253 -290
rect -253 -330 253 -324
<< properties >>
string FIXED_BBOX -258 -307 258 307
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.5 l 0.18 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc {+ 40} viadrn {- 40} viagate 100 viagb 100 viagr 0 viagl 0 viagt 0
<< end >>
