magic
tech sky130A
timestamp 1665556766
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_0
timestamp -19799
transform 1 0 -8 0 1 6
box -19 -24 249 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp -19799
transform 1 0 222 0 1 6
box -19 -24 65 296
<< end >>
