magic
tech sky130A
magscale 1 2
timestamp 1624218847
<< error_p >>
rect 198 51010 214 51026
rect 382 51010 398 51026
rect 182 50994 198 51010
rect 398 50994 414 51010
rect 61787 48353 61799 48356
rect 61746 48352 61799 48353
rect 61809 48352 61821 48356
rect 61859 48352 61871 48356
rect 61881 48352 61893 48356
rect 61746 48344 61788 48352
rect 61746 48327 61821 48344
rect 61822 48332 61833 48344
rect 61847 48332 61858 48344
rect 61738 48315 61746 48327
rect 61750 48310 61784 48327
rect 61787 48310 61821 48327
rect 61750 48231 61754 48265
rect 61780 48231 61784 48265
rect 61683 48194 61733 48196
rect 61700 48186 61722 48193
rect 61700 48185 61725 48186
rect 61733 48185 61735 48194
rect 61696 48178 61746 48185
rect 61696 48177 61742 48178
rect 61696 48173 61716 48177
rect 61708 48161 61716 48173
rect 61722 48161 61742 48177
rect 61708 48160 61742 48161
rect 61708 48153 61746 48160
rect 61722 48152 61725 48153
rect 61733 48144 61735 48153
rect 61750 48124 61753 48214
rect 61779 48183 61788 48211
rect 61777 48145 61788 48183
rect 61852 48173 61856 48327
rect 61859 48310 61864 48344
rect 61888 48313 61893 48344
rect 61894 48332 61905 48344
rect 62108 48327 62150 48353
rect 61882 48305 61954 48313
rect 61964 48305 62036 48313
rect 62040 48311 62044 48327
rect 62100 48319 62146 48327
rect 62100 48315 62116 48319
rect 62108 48312 62116 48315
rect 62142 48312 62146 48319
rect 62150 48315 62158 48327
rect 62096 48311 62162 48312
rect 61932 48275 61934 48291
rect 61904 48267 61934 48275
rect 61904 48263 61940 48267
rect 61904 48233 61912 48263
rect 61924 48233 61940 48263
rect 61932 48186 61934 48233
rect 62008 48206 62016 48275
rect 62040 48273 62050 48311
rect 62108 48303 62112 48311
rect 62162 48297 62212 48299
rect 62202 48293 62256 48297
rect 62202 48288 62222 48293
rect 62212 48273 62214 48288
rect 62044 48261 62050 48273
rect 61997 48196 62016 48206
rect 62008 48190 62016 48196
rect 62040 48227 62050 48261
rect 62108 48265 62112 48273
rect 62108 48231 62116 48265
rect 62142 48231 62146 48265
rect 62206 48263 62214 48273
rect 62222 48263 62223 48283
rect 62212 48247 62214 48263
rect 62233 48254 62236 48288
rect 62255 48263 62256 48283
rect 62265 48263 62272 48273
rect 62222 48247 62238 48253
rect 62240 48247 62256 48253
rect 62040 48199 62081 48227
rect 62040 48193 62059 48199
rect 61815 48139 61827 48173
rect 61837 48139 61857 48173
rect 61904 48152 61912 48186
rect 61924 48152 61940 48186
rect 61952 48180 61965 48186
rect 61986 48180 61999 48190
rect 61952 48156 61999 48180
rect 62008 48180 62029 48190
rect 62044 48183 62059 48193
rect 62008 48156 62037 48180
rect 62040 48165 62059 48183
rect 62069 48193 62083 48199
rect 62108 48193 62119 48231
rect 62270 48194 62320 48196
rect 62069 48165 62089 48193
rect 62108 48165 62117 48193
rect 62174 48185 62205 48193
rect 62273 48185 62304 48193
rect 62150 48178 62208 48185
rect 62174 48177 62208 48178
rect 62273 48177 62307 48185
rect 61952 48152 61965 48156
rect 61750 48073 61754 48107
rect 61780 48073 61784 48107
rect 61750 48026 61784 48030
rect 61750 48011 61754 48026
rect 61780 48011 61784 48026
rect 61746 47993 61788 48011
rect 61724 47987 61810 47993
rect 61852 47987 61856 48139
rect 61882 48115 61889 48143
rect 61932 48105 61934 48152
rect 62008 48143 62016 48156
rect 61986 48132 62013 48143
rect 62040 48115 62050 48165
rect 62108 48145 62112 48165
rect 62205 48161 62208 48177
rect 62304 48161 62307 48177
rect 62174 48160 62208 48161
rect 62150 48153 62208 48160
rect 62273 48153 62307 48161
rect 62320 48144 62322 48194
rect 61964 48105 62036 48113
rect 62044 48107 62050 48115
rect 62108 48107 62112 48115
rect 61904 48075 61912 48105
rect 61924 48075 61940 48105
rect 61904 48071 61940 48075
rect 61904 48063 61934 48071
rect 61932 48047 61934 48063
rect 62040 48035 62044 48103
rect 62108 48073 62116 48107
rect 62142 48073 62146 48107
rect 62162 48091 62212 48093
rect 62212 48075 62214 48091
rect 62222 48085 62238 48091
rect 62240 48085 62256 48091
rect 62233 48075 62256 48084
rect 62108 48065 62112 48073
rect 62206 48065 62214 48075
rect 62212 48041 62214 48065
rect 62222 48055 62223 48075
rect 62233 48050 62236 48075
rect 62255 48055 62256 48075
rect 62265 48065 62272 48075
rect 62222 48041 62256 48045
rect 62108 48035 62150 48036
rect 61882 48025 61954 48033
rect 62108 48028 62112 48035
rect 62003 47994 62008 48028
rect 62032 47994 62037 48028
rect 62075 48011 62146 48028
rect 62075 47994 62150 48011
rect 62108 47993 62150 47994
rect 62086 47987 62172 47993
rect 61746 47971 61788 47987
rect 62108 47971 62150 47987
rect 61683 47957 61733 47959
rect 61750 47957 61784 47971
rect 62112 47957 62146 47971
rect 62163 47957 62213 47959
rect 62265 47957 62315 47959
rect 61724 47949 61810 47957
rect 62086 47949 62172 47957
rect 61716 47915 61725 47949
rect 61726 47947 61759 47949
rect 61788 47947 61808 47949
rect 61726 47915 61808 47947
rect 62088 47947 62112 47949
rect 62137 47947 62146 47949
rect 62150 47947 62170 47949
rect 61724 47907 61810 47915
rect 61750 47891 61784 47907
rect 61724 47871 61746 47877
rect 61788 47871 61810 47877
rect 61852 47853 61856 47932
rect 62040 47877 62044 47932
rect 62088 47915 62170 47947
rect 62171 47915 62180 47949
rect 62188 47915 62205 47949
rect 62086 47907 62172 47915
rect 62213 47907 62215 47957
rect 62222 47915 62256 47949
rect 62273 47915 62290 47949
rect 62315 47907 62317 47957
rect 62112 47891 62146 47907
rect 62086 47871 62112 47877
rect 62150 47871 62172 47877
rect 62108 47853 62112 47871
rect 61746 47827 61788 47853
rect 62108 47827 62150 47853
rect 50984 398 51000 414
rect 51000 382 51016 398
rect 51000 198 51016 214
rect 50984 182 51000 198
use seal_ring_corner_abstract  seal_ring_corner_abstract_0 /usr/share/pdk/sky130A/libs.tech/magic/seal_ring_generator
timestamp 1624218757
transform 1 0 -200 0 1 -200
box 200 200 51216 51226
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_0 $PDKPATH/libs.ref/sky130_sram_macros/mag
timestamp 1624218757
transform 1 0 61708 0 1 47932
box -42 -105 650 424
<< labels >>
flabel space 251 52142 251 52142 0 FreeSans 9600 0 0 0 Unimplemented_rules
flabel space 62453 50878 62453 50878 0 FreeSans 9600 0 0 0 Unimplemented_rules
flabel space 137 53865 137 53865 0 FreeSans 9600 0 0 0 Exercise_8a
flabel space 62579 53228 62579 53228 0 FreeSans 9600 0 0 0 Exercise_8b
<< end >>
