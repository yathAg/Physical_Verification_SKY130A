magic
tech sky130A
magscale 1 2
timestamp 1626030382
<< metal3 >>
rect -3136 2872 3136 2900
rect -3136 -2872 3052 2872
rect 3116 -2872 3136 2872
rect -3136 -2900 3136 -2872
<< via3 >>
rect 3052 -2872 3116 2872
<< mimcap >>
rect -3036 2760 2964 2800
rect -3036 -2760 2332 2760
rect 2924 -2760 2964 2760
rect -3036 -2800 2964 -2760
<< mimcapcontact >>
rect 2332 -2760 2924 2760
<< metal4 >>
rect 3036 2872 3132 2888
rect 2331 2760 2925 2761
rect 2331 -2760 2332 2760
rect 2924 -2760 2925 2760
rect 2331 -2761 2925 -2760
rect 3036 -2872 3052 2872
rect 3116 -2872 3132 2872
rect 3036 -2888 3132 -2872
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX -3136 -2900 3064 2900
string parameters w 30.00 l 28.00 val 1.702k carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov -10
string library sky130
<< end >>
