magic
tech sky130A
magscale 1 2
timestamp 1624217268
<< checkpaint >>
rect 3491 -907 3859 -643
<< poly >>
rect 3491 -907 3859 -643
<< end >>
