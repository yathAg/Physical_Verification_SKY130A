magic
tech sky130A
magscale 1 2
timestamp 1624217737
<< metal2 >>
rect 4025 -872 4037 -805
rect 4104 -872 4128 -805
rect 4395 -872 4406 -805
<< via2 >>
rect 4037 -872 4104 -805
rect 4128 -872 4395 -805
<< metal3 >>
rect 4025 -805 4406 -800
rect 4025 -872 4037 -805
rect 4104 -872 4128 -805
rect 4395 -872 4406 -805
rect 4025 -877 4406 -872
<< end >>
