magic
tech sky130A
magscale 1 2
timestamp 1626030382
<< pwell >>
rect -5446 -2898 5446 2898
<< psubdiff >>
rect -5410 2828 -5314 2862
rect 5314 2828 5410 2862
rect -5410 2766 -5376 2828
rect 5376 2766 5410 2828
rect -5410 -2828 -5376 -2766
rect 5376 -2828 5410 -2766
rect -5410 -2862 -5314 -2828
rect 5314 -2862 5410 -2828
<< psubdiffcont >>
rect -5314 2828 5314 2862
rect -5410 -2766 -5376 2766
rect 5376 -2766 5410 2766
rect -5314 -2862 5314 -2828
<< xpolycontact >>
rect -5280 2300 -5142 2732
rect -5280 -2732 -5142 -2300
rect -4894 2300 -4756 2732
rect -4894 -2732 -4756 -2300
rect -4508 2300 -4370 2732
rect -4508 -2732 -4370 -2300
rect -4122 2300 -3984 2732
rect -4122 -2732 -3984 -2300
rect -3736 2300 -3598 2732
rect -3736 -2732 -3598 -2300
rect -3350 2300 -3212 2732
rect -3350 -2732 -3212 -2300
rect -2964 2300 -2826 2732
rect -2964 -2732 -2826 -2300
rect -2578 2300 -2440 2732
rect -2578 -2732 -2440 -2300
rect -2192 2300 -2054 2732
rect -2192 -2732 -2054 -2300
rect -1806 2300 -1668 2732
rect -1806 -2732 -1668 -2300
rect -1420 2300 -1282 2732
rect -1420 -2732 -1282 -2300
rect -1034 2300 -896 2732
rect -1034 -2732 -896 -2300
rect -648 2300 -510 2732
rect -648 -2732 -510 -2300
rect -262 2300 -124 2732
rect -262 -2732 -124 -2300
rect 124 2300 262 2732
rect 124 -2732 262 -2300
rect 510 2300 648 2732
rect 510 -2732 648 -2300
rect 896 2300 1034 2732
rect 896 -2732 1034 -2300
rect 1282 2300 1420 2732
rect 1282 -2732 1420 -2300
rect 1668 2300 1806 2732
rect 1668 -2732 1806 -2300
rect 2054 2300 2192 2732
rect 2054 -2732 2192 -2300
rect 2440 2300 2578 2732
rect 2440 -2732 2578 -2300
rect 2826 2300 2964 2732
rect 2826 -2732 2964 -2300
rect 3212 2300 3350 2732
rect 3212 -2732 3350 -2300
rect 3598 2300 3736 2732
rect 3598 -2732 3736 -2300
rect 3984 2300 4122 2732
rect 3984 -2732 4122 -2300
rect 4370 2300 4508 2732
rect 4370 -2732 4508 -2300
rect 4756 2300 4894 2732
rect 4756 -2732 4894 -2300
rect 5142 2300 5280 2732
rect 5142 -2732 5280 -2300
<< xpolyres >>
rect -5280 -2300 -5142 2300
rect -4894 -2300 -4756 2300
rect -4508 -2300 -4370 2300
rect -4122 -2300 -3984 2300
rect -3736 -2300 -3598 2300
rect -3350 -2300 -3212 2300
rect -2964 -2300 -2826 2300
rect -2578 -2300 -2440 2300
rect -2192 -2300 -2054 2300
rect -1806 -2300 -1668 2300
rect -1420 -2300 -1282 2300
rect -1034 -2300 -896 2300
rect -648 -2300 -510 2300
rect -262 -2300 -124 2300
rect 124 -2300 262 2300
rect 510 -2300 648 2300
rect 896 -2300 1034 2300
rect 1282 -2300 1420 2300
rect 1668 -2300 1806 2300
rect 2054 -2300 2192 2300
rect 2440 -2300 2578 2300
rect 2826 -2300 2964 2300
rect 3212 -2300 3350 2300
rect 3598 -2300 3736 2300
rect 3984 -2300 4122 2300
rect 4370 -2300 4508 2300
rect 4756 -2300 4894 2300
rect 5142 -2300 5280 2300
<< locali >>
rect -5410 2828 -5314 2862
rect 5314 2828 5410 2862
rect -5410 2766 -5376 2828
rect 5376 2766 5410 2828
rect -5410 -2828 -5376 -2766
rect 5376 -2828 5410 -2766
rect -5410 -2862 -5314 -2828
rect 5314 -2862 5410 -2828
<< viali >>
rect -5410 -2545 -5376 2545
rect 5376 -2545 5410 2545
rect -4838 -2862 4838 -2828
<< metal1 >>
rect -5416 2545 -5370 2557
rect -5416 -2545 -5410 2545
rect -5376 -2545 -5370 2545
rect -5416 -2557 -5370 -2545
rect 5370 2545 5416 2557
rect 5370 -2545 5376 2545
rect 5410 -2545 5416 2545
rect 5370 -2557 5416 -2545
rect -4850 -2828 4850 -2822
rect -4850 -2862 -4838 -2828
rect 4838 -2862 4850 -2828
rect -4850 -2868 4850 -2862
<< res0p69 >>
rect -5282 -2302 -5140 2302
rect -4896 -2302 -4754 2302
rect -4510 -2302 -4368 2302
rect -4124 -2302 -3982 2302
rect -3738 -2302 -3596 2302
rect -3352 -2302 -3210 2302
rect -2966 -2302 -2824 2302
rect -2580 -2302 -2438 2302
rect -2194 -2302 -2052 2302
rect -1808 -2302 -1666 2302
rect -1422 -2302 -1280 2302
rect -1036 -2302 -894 2302
rect -650 -2302 -508 2302
rect -264 -2302 -122 2302
rect 122 -2302 264 2302
rect 508 -2302 650 2302
rect 894 -2302 1036 2302
rect 1280 -2302 1422 2302
rect 1666 -2302 1808 2302
rect 2052 -2302 2194 2302
rect 2438 -2302 2580 2302
rect 2824 -2302 2966 2302
rect 3210 -2302 3352 2302
rect 3596 -2302 3738 2302
rect 3982 -2302 4124 2302
rect 4368 -2302 4510 2302
rect 4754 -2302 4896 2302
rect 5140 -2302 5282 2302
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p69
string FIXED_BBOX -5393 -2845 5393 2845
string parameters w 0.69 l 23.0 m 1 nx 28 wmin 0.690 lmin 0.50 rho 2000 val 66.722k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 wmax 0.690 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 0 viagb 90 viagt 0 viagl 90 viagr 90
string library sky130
<< end >>
