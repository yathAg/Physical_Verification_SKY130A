magic
tech sky130A
magscale 1 2
timestamp 1626025383
<< locali >>
rect 5733 12087 5767 12257
rect 7573 10523 7607 10625
rect 9321 10591 9355 10761
rect 2697 8959 2731 9129
rect 9965 9027 9999 9129
rect 11069 9027 11103 9129
rect 9137 8347 9171 8449
rect 5457 7735 5491 8041
rect 6009 6715 6043 6817
rect 10333 6307 10367 6409
rect 9505 5559 9539 5729
rect 5825 4607 5859 4777
rect 6653 4675 6687 4777
rect 7481 3145 7573 3179
rect 5181 2975 5215 3145
rect 7481 2975 7515 3145
rect 11437 2975 11471 3145
rect 6377 2295 6411 2397
rect 10517 2363 10551 2601
rect 9045 1751 9079 1921
rect 11529 1887 11563 1989
rect 11713 1411 11747 1513
<< viali >>
rect 4905 15657 4939 15691
rect 4813 15589 4847 15623
rect 4169 15521 4203 15555
rect 5641 15521 5675 15555
rect 6193 15521 6227 15555
rect 6837 15521 6871 15555
rect 7481 15521 7515 15555
rect 9413 15521 9447 15555
rect 10241 15521 10275 15555
rect 5089 15453 5123 15487
rect 8033 15453 8067 15487
rect 8585 15453 8619 15487
rect 6101 15385 6135 15419
rect 8493 15385 8527 15419
rect 9229 15385 9263 15419
rect 4077 15317 4111 15351
rect 4445 15317 4479 15351
rect 5457 15317 5491 15351
rect 6653 15317 6687 15351
rect 7297 15317 7331 15351
rect 10149 15317 10183 15351
rect 6009 15113 6043 15147
rect 10609 15045 10643 15079
rect 7205 14977 7239 15011
rect 7389 14977 7423 15011
rect 9873 14977 9907 15011
rect 10057 14977 10091 15011
rect 11161 14977 11195 15011
rect 3801 14909 3835 14943
rect 4721 14909 4755 14943
rect 6009 14909 6043 14943
rect 7849 14909 7883 14943
rect 11069 14909 11103 14943
rect 4537 14841 4571 14875
rect 8585 14841 8619 14875
rect 8769 14841 8803 14875
rect 6745 14773 6779 14807
rect 7113 14773 7147 14807
rect 9413 14773 9447 14807
rect 9781 14773 9815 14807
rect 10977 14773 11011 14807
rect 2237 14569 2271 14603
rect 11069 14569 11103 14603
rect 3893 14501 3927 14535
rect 5181 14501 5215 14535
rect 5273 14501 5307 14535
rect 7389 14501 7423 14535
rect 2145 14433 2179 14467
rect 3157 14433 3191 14467
rect 4721 14433 4755 14467
rect 5549 14433 5583 14467
rect 6469 14433 6503 14467
rect 7481 14433 7515 14467
rect 8217 14433 8251 14467
rect 9229 14433 9263 14467
rect 10701 14433 10735 14467
rect 11713 14433 11747 14467
rect 2329 14365 2363 14399
rect 4445 14365 4479 14399
rect 7941 14365 7975 14399
rect 8769 14365 8803 14399
rect 11161 14365 11195 14399
rect 2973 14297 3007 14331
rect 3985 14297 4019 14331
rect 6837 14297 6871 14331
rect 8677 14297 8711 14331
rect 10517 14297 10551 14331
rect 1777 14229 1811 14263
rect 11529 14229 11563 14263
rect 5917 14025 5951 14059
rect 6929 13957 6963 13991
rect 9045 13957 9079 13991
rect 9965 13957 9999 13991
rect 10793 13957 10827 13991
rect 12265 13957 12299 13991
rect 4905 13889 4939 13923
rect 5365 13889 5399 13923
rect 5457 13889 5491 13923
rect 6469 13889 6503 13923
rect 7021 13889 7055 13923
rect 9505 13889 9539 13923
rect 10057 13889 10091 13923
rect 10885 13889 10919 13923
rect 1869 13821 1903 13855
rect 3341 13821 3375 13855
rect 4813 13821 4847 13855
rect 7573 13821 7607 13855
rect 8769 13821 8803 13855
rect 10333 13821 10367 13855
rect 11713 13821 11747 13855
rect 12449 13821 12483 13855
rect 13185 13821 13219 13855
rect 2513 13753 2547 13787
rect 2789 13753 2823 13787
rect 11897 13753 11931 13787
rect 5549 13685 5583 13719
rect 11253 13685 11287 13719
rect 11345 13685 11379 13719
rect 13001 13685 13035 13719
rect 2881 13481 2915 13515
rect 3893 13481 3927 13515
rect 1685 13413 1719 13447
rect 2421 13413 2455 13447
rect 4629 13413 4663 13447
rect 5181 13413 5215 13447
rect 6837 13413 6871 13447
rect 8493 13413 8527 13447
rect 8677 13413 8711 13447
rect 10241 13413 10275 13447
rect 10517 13413 10551 13447
rect 11989 13413 12023 13447
rect 1961 13345 1995 13379
rect 2973 13345 3007 13379
rect 3525 13345 3559 13379
rect 4077 13345 4111 13379
rect 4445 13345 4479 13379
rect 5365 13345 5399 13379
rect 5825 13345 5859 13379
rect 6009 13345 6043 13379
rect 6653 13345 6687 13379
rect 7573 13345 7607 13379
rect 8033 13345 8067 13379
rect 9137 13345 9171 13379
rect 9597 13345 9631 13379
rect 11069 13345 11103 13379
rect 11713 13345 11747 13379
rect 12725 13345 12759 13379
rect 12909 13345 12943 13379
rect 13369 13345 13403 13379
rect 2513 13277 2547 13311
rect 7849 13277 7883 13311
rect 3341 13209 3375 13243
rect 1593 13141 1627 13175
rect 5089 13141 5123 13175
rect 5733 13141 5767 13175
rect 9229 13141 9263 13175
rect 13185 13141 13219 13175
rect 5917 12937 5951 12971
rect 8217 12937 8251 12971
rect 9781 12937 9815 12971
rect 2881 12869 2915 12903
rect 9505 12869 9539 12903
rect 1593 12801 1627 12835
rect 2973 12801 3007 12835
rect 3985 12801 4019 12835
rect 5365 12801 5399 12835
rect 6837 12801 6871 12835
rect 8861 12801 8895 12835
rect 9045 12801 9079 12835
rect 10241 12801 10275 12835
rect 10425 12801 10459 12835
rect 11345 12801 11379 12835
rect 1777 12733 1811 12767
rect 2421 12733 2455 12767
rect 3525 12733 3559 12767
rect 4537 12733 4571 12767
rect 5549 12733 5583 12767
rect 7665 12733 7699 12767
rect 8309 12733 8343 12767
rect 10149 12733 10183 12767
rect 10793 12733 10827 12767
rect 11713 12733 11747 12767
rect 13185 12733 13219 12767
rect 4077 12665 4111 12699
rect 4721 12665 4755 12699
rect 4905 12665 4939 12699
rect 5457 12665 5491 12699
rect 6929 12665 6963 12699
rect 8493 12665 8527 12699
rect 11253 12665 11287 12699
rect 13277 12665 13311 12699
rect 1685 12597 1719 12631
rect 2145 12597 2179 12631
rect 7021 12597 7055 12631
rect 7389 12597 7423 12631
rect 7757 12597 7791 12631
rect 9137 12597 9171 12631
rect 4353 12393 4387 12427
rect 5917 12393 5951 12427
rect 7297 12393 7331 12427
rect 9321 12393 9355 12427
rect 9781 12393 9815 12427
rect 12357 12393 12391 12427
rect 13093 12393 13127 12427
rect 3065 12325 3099 12359
rect 11713 12325 11747 12359
rect 1501 12257 1535 12291
rect 2789 12257 2823 12291
rect 3341 12257 3375 12291
rect 4261 12257 4295 12291
rect 4905 12257 4939 12291
rect 5181 12257 5215 12291
rect 5457 12257 5491 12291
rect 5733 12257 5767 12291
rect 6101 12257 6135 12291
rect 6377 12257 6411 12291
rect 6745 12257 6779 12291
rect 7481 12257 7515 12291
rect 7757 12257 7791 12291
rect 7941 12257 7975 12291
rect 8493 12257 8527 12291
rect 8677 12257 8711 12291
rect 9689 12257 9723 12291
rect 10333 12257 10367 12291
rect 10517 12257 10551 12291
rect 11161 12257 11195 12291
rect 11621 12257 11655 12291
rect 13185 12257 13219 12291
rect 4537 12189 4571 12223
rect 5365 12189 5399 12223
rect 3893 12121 3927 12155
rect 5277 12121 5311 12155
rect 7665 12189 7699 12223
rect 9965 12189 9999 12223
rect 12449 12189 12483 12223
rect 12541 12189 12575 12223
rect 6197 12121 6231 12155
rect 6285 12121 6319 12155
rect 7573 12121 7607 12155
rect 3525 12053 3559 12087
rect 5733 12053 5767 12087
rect 6837 12053 6871 12087
rect 8309 12053 8343 12087
rect 8493 12053 8527 12087
rect 10609 12053 10643 12087
rect 11989 12053 12023 12087
rect 6009 11849 6043 11883
rect 6561 11849 6595 11883
rect 11713 11849 11747 11883
rect 5089 11781 5123 11815
rect 6929 11781 6963 11815
rect 8309 11781 8343 11815
rect 9501 11781 9535 11815
rect 10885 11781 10919 11815
rect 13185 11781 13219 11815
rect 2237 11713 2271 11747
rect 2329 11713 2363 11747
rect 7021 11713 7055 11747
rect 7113 11713 7147 11747
rect 8401 11713 8435 11747
rect 9413 11713 9447 11747
rect 10517 11713 10551 11747
rect 12357 11713 12391 11747
rect 13277 11713 13311 11747
rect 3157 11645 3191 11679
rect 3433 11645 3467 11679
rect 4169 11645 4203 11679
rect 5917 11645 5951 11679
rect 6837 11645 6871 11679
rect 7205 11645 7239 11679
rect 8033 11645 8067 11679
rect 8217 11645 8251 11679
rect 8493 11645 8527 11679
rect 8677 11645 8711 11679
rect 9321 11645 9355 11679
rect 9597 11645 9631 11679
rect 9873 11645 9907 11679
rect 10977 11645 11011 11679
rect 11161 11645 11195 11679
rect 12725 11645 12759 11679
rect 2145 11577 2179 11611
rect 2789 11577 2823 11611
rect 2973 11577 3007 11611
rect 4353 11577 4387 11611
rect 5273 11577 5307 11611
rect 5641 11577 5675 11611
rect 10149 11577 10183 11611
rect 10333 11577 10367 11611
rect 12081 11577 12115 11611
rect 1777 11509 1811 11543
rect 4629 11509 4663 11543
rect 5365 11509 5399 11543
rect 5457 11509 5491 11543
rect 12173 11509 12207 11543
rect 7665 11305 7699 11339
rect 8033 11305 8067 11339
rect 9597 11305 9631 11339
rect 11069 11305 11103 11339
rect 3893 11237 3927 11271
rect 3985 11237 4019 11271
rect 5641 11237 5675 11271
rect 6101 11237 6135 11271
rect 8125 11237 8159 11271
rect 10977 11237 11011 11271
rect 13369 11237 13403 11271
rect 1777 11169 1811 11203
rect 2421 11169 2455 11203
rect 2697 11169 2731 11203
rect 3525 11169 3559 11203
rect 4445 11169 4479 11203
rect 4905 11169 4939 11203
rect 5181 11169 5215 11203
rect 5457 11169 5491 11203
rect 6009 11169 6043 11203
rect 6469 11169 6503 11203
rect 6745 11169 6779 11203
rect 7021 11169 7055 11203
rect 7205 11169 7239 11203
rect 9873 11169 9907 11203
rect 9965 11169 9999 11203
rect 10333 11169 10367 11203
rect 11805 11169 11839 11203
rect 13277 11169 13311 11203
rect 2973 11101 3007 11135
rect 5273 11101 5307 11135
rect 6929 11101 6963 11135
rect 8217 11101 8251 11135
rect 11161 11101 11195 11135
rect 3065 11033 3099 11067
rect 4721 11033 4755 11067
rect 6837 11033 6871 11067
rect 10057 10965 10091 10999
rect 10149 10965 10183 10999
rect 10609 10965 10643 10999
rect 2881 10761 2915 10795
rect 6837 10761 6871 10795
rect 8677 10761 8711 10795
rect 9321 10761 9355 10795
rect 9689 10761 9723 10795
rect 11805 10761 11839 10795
rect 4629 10693 4663 10727
rect 5917 10693 5951 10727
rect 5549 10625 5583 10659
rect 7021 10625 7055 10659
rect 7573 10625 7607 10659
rect 1593 10557 1627 10591
rect 1869 10557 1903 10591
rect 2329 10557 2363 10591
rect 2697 10557 2731 10591
rect 3157 10557 3191 10591
rect 4169 10557 4203 10591
rect 5457 10557 5491 10591
rect 5641 10557 5675 10591
rect 5733 10557 5767 10591
rect 7113 10557 7147 10591
rect 10885 10625 10919 10659
rect 7665 10557 7699 10591
rect 8677 10557 8711 10591
rect 8861 10557 8895 10591
rect 9321 10557 9355 10591
rect 9413 10557 9447 10591
rect 10057 10557 10091 10591
rect 10425 10557 10459 10591
rect 11069 10557 11103 10591
rect 11713 10557 11747 10591
rect 11897 10557 11931 10591
rect 12357 10557 12391 10591
rect 13001 10557 13035 10591
rect 13277 10557 13311 10591
rect 1501 10489 1535 10523
rect 2421 10489 2455 10523
rect 6837 10489 6871 10523
rect 7573 10489 7607 10523
rect 7849 10489 7883 10523
rect 8033 10489 8067 10523
rect 9597 10489 9631 10523
rect 10609 10489 10643 10523
rect 7297 10421 7331 10455
rect 9045 10421 9079 10455
rect 10241 10421 10275 10455
rect 10333 10421 10367 10455
rect 11253 10421 11287 10455
rect 10057 10217 10091 10251
rect 2973 10149 3007 10183
rect 9229 10149 9263 10183
rect 13093 10149 13127 10183
rect 1409 10081 1443 10115
rect 2697 10081 2731 10115
rect 3341 10081 3375 10115
rect 3985 10081 4019 10115
rect 4261 10081 4295 10115
rect 5181 10081 5215 10115
rect 5457 10081 5491 10115
rect 5549 10081 5583 10115
rect 6561 10081 6595 10115
rect 6745 10081 6779 10115
rect 6929 10081 6963 10115
rect 7573 10081 7607 10115
rect 7849 10081 7883 10115
rect 8033 10081 8067 10115
rect 8309 10081 8343 10115
rect 8585 10081 8619 10115
rect 9137 10081 9171 10115
rect 9321 10081 9355 10115
rect 9505 10081 9539 10115
rect 9965 10081 9999 10115
rect 10425 10081 10459 10115
rect 13001 10081 13035 10115
rect 5273 10013 5307 10047
rect 7389 10013 7423 10047
rect 10701 10013 10735 10047
rect 12541 10013 12575 10047
rect 3985 9945 4019 9979
rect 6285 9945 6319 9979
rect 7665 9945 7699 9979
rect 7757 9945 7791 9979
rect 8585 9945 8619 9979
rect 3525 9877 3559 9911
rect 4905 9877 4939 9911
rect 5365 9877 5399 9911
rect 6653 9877 6687 9911
rect 6837 9877 6871 9911
rect 12173 9877 12207 9911
rect 1409 9673 1443 9707
rect 3341 9673 3375 9707
rect 5549 9673 5583 9707
rect 5733 9673 5767 9707
rect 7113 9673 7147 9707
rect 10793 9673 10827 9707
rect 12265 9673 12299 9707
rect 8953 9605 8987 9639
rect 9873 9605 9907 9639
rect 2053 9537 2087 9571
rect 6653 9537 6687 9571
rect 8289 9537 8323 9571
rect 9781 9537 9815 9571
rect 11253 9537 11287 9571
rect 11805 9537 11839 9571
rect 12817 9537 12851 9571
rect 1777 9469 1811 9503
rect 2789 9469 2823 9503
rect 3249 9469 3283 9503
rect 3525 9469 3559 9503
rect 4629 9469 4663 9503
rect 6745 9469 6779 9503
rect 8585 9469 8619 9503
rect 9085 9469 9119 9503
rect 9228 9469 9262 9503
rect 9505 9469 9539 9503
rect 10057 9469 10091 9503
rect 10149 9469 10183 9503
rect 11069 9469 11103 9503
rect 11897 9469 11931 9503
rect 12633 9469 12667 9503
rect 3985 9401 4019 9435
rect 5733 9401 5767 9435
rect 5917 9401 5951 9435
rect 7205 9401 7239 9435
rect 7389 9401 7423 9435
rect 7849 9401 7883 9435
rect 8033 9401 8067 9435
rect 8493 9401 8527 9435
rect 9321 9401 9355 9435
rect 10701 9401 10735 9435
rect 1869 9333 1903 9367
rect 2881 9333 2915 9367
rect 8401 9333 8435 9367
rect 10333 9333 10367 9367
rect 12725 9333 12759 9367
rect 1961 9129 1995 9163
rect 2697 9129 2731 9163
rect 4261 9129 4295 9163
rect 9965 9129 9999 9163
rect 10793 9129 10827 9163
rect 11069 9129 11103 9163
rect 12725 9129 12759 9163
rect 1593 9061 1627 9095
rect 1869 8993 1903 9027
rect 2329 8993 2363 9027
rect 7113 9061 7147 9095
rect 10425 9061 10459 9095
rect 10517 9061 10551 9095
rect 11897 9061 11931 9095
rect 3893 8993 3927 9027
rect 4261 8993 4295 9027
rect 4905 8993 4939 9027
rect 4997 8993 5031 9027
rect 5181 8993 5215 9027
rect 7849 8993 7883 9027
rect 8033 8993 8067 9027
rect 8309 8993 8343 9027
rect 9137 8993 9171 9027
rect 9321 8993 9355 9027
rect 9505 8993 9539 9027
rect 9965 8993 9999 9027
rect 10149 8993 10183 9027
rect 10297 8993 10331 9027
rect 10614 8993 10648 9027
rect 11069 8993 11103 9027
rect 11161 8993 11195 9027
rect 11345 8993 11379 9027
rect 11805 8993 11839 9027
rect 12265 8993 12299 9027
rect 12909 8993 12943 9027
rect 13369 8993 13403 9027
rect 2697 8925 2731 8959
rect 2789 8925 2823 8959
rect 3341 8925 3375 8959
rect 5641 8925 5675 8959
rect 7389 8925 7423 8959
rect 8125 8925 8159 8959
rect 8217 8925 8251 8959
rect 9413 8925 9447 8959
rect 9598 8925 9632 8959
rect 12357 8925 12391 8959
rect 1501 8857 1535 8891
rect 2513 8857 2547 8891
rect 2881 8857 2915 8891
rect 5089 8857 5123 8891
rect 8493 8857 8527 8891
rect 13185 8857 13219 8891
rect 4721 8789 4755 8823
rect 9781 8789 9815 8823
rect 11253 8789 11287 8823
rect 5365 8585 5399 8619
rect 6101 8585 6135 8619
rect 7113 8585 7147 8619
rect 8677 8585 8711 8619
rect 6929 8517 6963 8551
rect 8217 8517 8251 8551
rect 10517 8517 10551 8551
rect 13093 8517 13127 8551
rect 2053 8449 2087 8483
rect 7021 8449 7055 8483
rect 9137 8449 9171 8483
rect 9321 8449 9355 8483
rect 12725 8449 12759 8483
rect 1777 8381 1811 8415
rect 2697 8381 2731 8415
rect 3341 8381 3375 8415
rect 3617 8381 3651 8415
rect 5917 8381 5951 8415
rect 6837 8381 6871 8415
rect 7205 8381 7239 8415
rect 7665 8381 7699 8415
rect 8038 8381 8072 8415
rect 8769 8381 8803 8415
rect 8953 8381 8987 8415
rect 9229 8381 9263 8415
rect 9505 8381 9539 8415
rect 9597 8381 9631 8415
rect 9781 8381 9815 8415
rect 10333 8381 10367 8415
rect 10517 8381 10551 8415
rect 10977 8381 11011 8415
rect 12449 8381 12483 8415
rect 13277 8381 13311 8415
rect 1869 8313 1903 8347
rect 2421 8313 2455 8347
rect 3893 8313 3927 8347
rect 7849 8313 7883 8347
rect 7941 8313 7975 8347
rect 9137 8313 9171 8347
rect 10149 8313 10183 8347
rect 11069 8313 11103 8347
rect 1409 8245 1443 8279
rect 6561 8245 6595 8279
rect 12081 8245 12115 8279
rect 12541 8245 12575 8279
rect 4721 8041 4755 8075
rect 4905 8041 4939 8075
rect 5457 8041 5491 8075
rect 5641 8041 5675 8075
rect 6193 8041 6227 8075
rect 6561 8041 6595 8075
rect 9781 8041 9815 8075
rect 11989 8041 12023 8075
rect 4077 7973 4111 8007
rect 1501 7905 1535 7939
rect 2973 7905 3007 7939
rect 3341 7905 3375 7939
rect 4903 7905 4937 7939
rect 5365 7905 5399 7939
rect 3893 7837 3927 7871
rect 2973 7769 3007 7803
rect 3525 7769 3559 7803
rect 7941 7973 7975 8007
rect 9413 7973 9447 8007
rect 9505 7973 9539 8007
rect 10517 7973 10551 8007
rect 13093 7973 13127 8007
rect 5825 7905 5859 7939
rect 6653 7905 6687 7939
rect 7205 7905 7239 7939
rect 8033 7905 8067 7939
rect 9137 7905 9171 7939
rect 9285 7905 9319 7939
rect 9643 7905 9677 7939
rect 12357 7905 12391 7939
rect 13277 7905 13311 7939
rect 6837 7837 6871 7871
rect 7849 7837 7883 7871
rect 10241 7837 10275 7871
rect 5273 7701 5307 7735
rect 5457 7701 5491 7735
rect 7297 7701 7331 7735
rect 8401 7701 8435 7735
rect 10149 7497 10183 7531
rect 13001 7497 13035 7531
rect 5365 7429 5399 7463
rect 9505 7429 9539 7463
rect 12541 7429 12575 7463
rect 1961 7361 1995 7395
rect 2513 7361 2547 7395
rect 5273 7361 5307 7395
rect 7021 7361 7055 7395
rect 8016 7361 8050 7395
rect 8309 7361 8343 7395
rect 10793 7361 10827 7395
rect 11345 7361 11379 7395
rect 12633 7361 12667 7395
rect 1501 7293 1535 7327
rect 2421 7293 2455 7327
rect 2973 7293 3007 7327
rect 3433 7293 3467 7327
rect 3893 7293 3927 7327
rect 5825 7293 5859 7327
rect 6837 7293 6871 7327
rect 7757 7293 7791 7327
rect 8094 7293 8128 7327
rect 9229 7293 9263 7327
rect 9321 7293 9355 7327
rect 9597 7293 9631 7327
rect 10149 7293 10183 7327
rect 10333 7293 10367 7327
rect 12081 7293 12115 7327
rect 12909 7293 12943 7327
rect 2789 7225 2823 7259
rect 4537 7225 4571 7259
rect 4813 7225 4847 7259
rect 7573 7225 7607 7259
rect 11253 7225 11287 7259
rect 1685 7157 1719 7191
rect 3617 7157 3651 7191
rect 6469 7157 6503 7191
rect 6929 7157 6963 7191
rect 8217 7157 8251 7191
rect 9045 7157 9079 7191
rect 9965 7157 9999 7191
rect 3157 6953 3191 6987
rect 2513 6885 2547 6919
rect 8493 6885 8527 6919
rect 11253 6885 11287 6919
rect 1593 6817 1627 6851
rect 2237 6817 2271 6851
rect 3065 6817 3099 6851
rect 3893 6817 3927 6851
rect 4353 6817 4387 6851
rect 5825 6817 5859 6851
rect 6009 6817 6043 6851
rect 8033 6817 8067 6851
rect 8309 6817 8343 6851
rect 9137 6817 9171 6851
rect 9689 6817 9723 6851
rect 11161 6817 11195 6851
rect 2652 6750 2686 6784
rect 2973 6749 3007 6783
rect 13093 6749 13127 6783
rect 13369 6749 13403 6783
rect 4077 6681 4111 6715
rect 5825 6681 5859 6715
rect 6009 6681 6043 6715
rect 3525 6613 3559 6647
rect 6285 6613 6319 6647
rect 7769 6613 7803 6647
rect 8585 6613 8619 6647
rect 9229 6613 9263 6647
rect 11621 6613 11655 6647
rect 7021 6409 7055 6443
rect 10333 6409 10367 6443
rect 1869 6341 1903 6375
rect 2513 6341 2547 6375
rect 4537 6341 4571 6375
rect 7389 6341 7423 6375
rect 9045 6341 9079 6375
rect 11069 6341 11103 6375
rect 1409 6273 1443 6307
rect 1961 6273 1995 6307
rect 5273 6273 5307 6307
rect 5457 6273 5491 6307
rect 10333 6273 10367 6307
rect 11989 6273 12023 6307
rect 2513 6205 2547 6239
rect 3801 6205 3835 6239
rect 4353 6205 4387 6239
rect 5181 6205 5215 6239
rect 6101 6205 6135 6239
rect 6929 6205 6963 6239
rect 7113 6205 7147 6239
rect 7631 6205 7665 6239
rect 7757 6205 7791 6239
rect 7849 6205 7883 6239
rect 8033 6205 8067 6239
rect 8585 6205 8619 6239
rect 8861 6205 8895 6239
rect 8953 6205 8987 6239
rect 9137 6205 9171 6239
rect 9735 6205 9769 6239
rect 9873 6205 9907 6239
rect 10149 6205 10183 6239
rect 10517 6205 10551 6239
rect 10890 6205 10924 6239
rect 12449 6205 12483 6239
rect 12909 6205 12943 6239
rect 13369 6205 13403 6239
rect 6009 6137 6043 6171
rect 10241 6137 10275 6171
rect 10701 6137 10735 6171
rect 10793 6137 10827 6171
rect 11805 6137 11839 6171
rect 4813 6069 4847 6103
rect 9597 6069 9631 6103
rect 12265 6069 12299 6103
rect 12725 6069 12759 6103
rect 13185 6069 13219 6103
rect 1409 5865 1443 5899
rect 1869 5865 1903 5899
rect 5273 5865 5307 5899
rect 10977 5865 11011 5899
rect 2789 5797 2823 5831
rect 4629 5797 4663 5831
rect 9229 5797 9263 5831
rect 11069 5797 11103 5831
rect 11713 5797 11747 5831
rect 1777 5729 1811 5763
rect 3341 5729 3375 5763
rect 4077 5729 4111 5763
rect 4537 5729 4571 5763
rect 5365 5729 5399 5763
rect 5641 5729 5675 5763
rect 8217 5729 8251 5763
rect 8309 5729 8343 5763
rect 8585 5729 8619 5763
rect 9137 5729 9171 5763
rect 9505 5729 9539 5763
rect 9597 5729 9631 5763
rect 9873 5729 9907 5763
rect 10149 5729 10183 5763
rect 10333 5729 10367 5763
rect 2053 5661 2087 5695
rect 2881 5661 2915 5695
rect 9965 5661 9999 5695
rect 11437 5661 11471 5695
rect 5898 5525 5932 5559
rect 7389 5525 7423 5559
rect 8033 5525 8067 5559
rect 8493 5525 8527 5559
rect 9505 5525 9539 5559
rect 13185 5525 13219 5559
rect 8769 5321 8803 5355
rect 11253 5321 11287 5355
rect 12541 5253 12575 5287
rect 7297 5185 7331 5219
rect 9505 5185 9539 5219
rect 9781 5185 9815 5219
rect 12705 5185 12739 5219
rect 13185 5185 13219 5219
rect 1593 5117 1627 5151
rect 3893 5117 3927 5151
rect 6009 5117 6043 5151
rect 6469 5117 6503 5151
rect 11897 5117 11931 5151
rect 12817 5117 12851 5151
rect 3617 5049 3651 5083
rect 5733 5049 5767 5083
rect 13093 5049 13127 5083
rect 1777 4981 1811 5015
rect 2145 4981 2179 5015
rect 4261 4981 4295 5015
rect 6561 4981 6595 5015
rect 11805 4981 11839 5015
rect 3968 4777 4002 4811
rect 5273 4777 5307 4811
rect 5825 4777 5859 4811
rect 4261 4709 4295 4743
rect 1593 4641 1627 4675
rect 2053 4641 2087 4675
rect 2421 4641 2455 4675
rect 2697 4641 2731 4675
rect 3341 4641 3375 4675
rect 3525 4641 3559 4675
rect 4164 4641 4198 4675
rect 4353 4641 4387 4675
rect 4537 4641 4571 4675
rect 4997 4641 5031 4675
rect 6653 4777 6687 4811
rect 13277 4777 13311 4811
rect 6285 4709 6319 4743
rect 9137 4709 9171 4743
rect 6141 4641 6175 4675
rect 6377 4641 6411 4675
rect 6561 4641 6595 4675
rect 6653 4641 6687 4675
rect 6837 4641 6871 4675
rect 7297 4641 7331 4675
rect 8033 4641 8067 4675
rect 8309 4641 8343 4675
rect 8493 4641 8527 4675
rect 9321 4641 9355 4675
rect 9690 4641 9724 4675
rect 9873 4641 9907 4675
rect 10517 4641 10551 4675
rect 10977 4641 11011 4675
rect 11529 4641 11563 4675
rect 2329 4573 2363 4607
rect 2973 4573 3007 4607
rect 4813 4573 4847 4607
rect 5365 4573 5399 4607
rect 5825 4573 5859 4607
rect 6929 4573 6963 4607
rect 9505 4573 9539 4607
rect 9597 4573 9631 4607
rect 10149 4573 10183 4607
rect 10701 4573 10735 4607
rect 11805 4573 11839 4607
rect 1501 4505 1535 4539
rect 3065 4505 3099 4539
rect 6009 4505 6043 4539
rect 7941 4505 7975 4539
rect 8677 4505 8711 4539
rect 10241 4505 10275 4539
rect 1961 4437 1995 4471
rect 7389 4437 7423 4471
rect 8493 4437 8527 4471
rect 11069 4437 11103 4471
rect 3065 4233 3099 4267
rect 9768 4233 9802 4267
rect 11805 4233 11839 4267
rect 8125 4097 8159 4131
rect 8217 4097 8251 4131
rect 9137 4097 9171 4131
rect 11253 4097 11287 4131
rect 1777 4029 1811 4063
rect 1961 4029 1995 4063
rect 2053 4029 2087 4063
rect 2146 4029 2180 4063
rect 2973 4029 3007 4063
rect 3495 4029 3529 4063
rect 5917 4029 5951 4063
rect 6740 4029 6774 4063
rect 7113 4029 7147 4063
rect 7941 4029 7975 4063
rect 8345 4029 8379 4063
rect 8493 4029 8527 4063
rect 9505 4029 9539 4063
rect 11937 4029 11971 4063
rect 12173 4029 12207 4063
rect 12357 4029 12391 4063
rect 12633 4029 12667 4063
rect 13277 4029 13311 4063
rect 2421 3961 2455 3995
rect 5641 3961 5675 3995
rect 6837 3961 6871 3995
rect 6929 3961 6963 3995
rect 8769 3961 8803 3995
rect 8953 3961 8987 3995
rect 12081 3961 12115 3995
rect 3433 3893 3467 3927
rect 3617 3893 3651 3927
rect 4169 3893 4203 3927
rect 6553 3893 6587 3927
rect 7849 3893 7883 3927
rect 12725 3893 12759 3927
rect 13093 3893 13127 3927
rect 2605 3689 2639 3723
rect 5365 3689 5399 3723
rect 5457 3689 5491 3723
rect 5641 3689 5675 3723
rect 10517 3689 10551 3723
rect 3157 3621 3191 3655
rect 1501 3553 1535 3587
rect 1685 3553 1719 3587
rect 1961 3553 1995 3587
rect 2237 3553 2271 3587
rect 2881 3553 2915 3587
rect 3249 3553 3283 3587
rect 4261 3553 4295 3587
rect 4537 3553 4571 3587
rect 5181 3553 5215 3587
rect 5549 3553 5583 3587
rect 6285 3553 6319 3587
rect 6469 3553 6503 3587
rect 6929 3553 6963 3587
rect 7113 3553 7147 3587
rect 7481 3553 7515 3587
rect 7941 3553 7975 3587
rect 8217 3553 8251 3587
rect 8401 3553 8435 3587
rect 8585 3553 8619 3587
rect 9137 3553 9171 3587
rect 9321 3553 9355 3587
rect 9689 3553 9723 3587
rect 9965 3553 9999 3587
rect 10149 3553 10183 3587
rect 10609 3553 10643 3587
rect 10793 3553 10827 3587
rect 10978 3553 11012 3587
rect 11161 3553 11195 3587
rect 2769 3485 2803 3519
rect 4149 3485 4183 3519
rect 4629 3485 4663 3519
rect 7757 3485 7791 3519
rect 7849 3485 7883 3519
rect 9229 3485 9263 3519
rect 10885 3485 10919 3519
rect 11529 3485 11563 3519
rect 11805 3485 11839 3519
rect 13277 3485 13311 3519
rect 1869 3417 1903 3451
rect 3985 3417 4019 3451
rect 6101 3349 6135 3383
rect 6469 3349 6503 3383
rect 4445 3145 4479 3179
rect 5181 3145 5215 3179
rect 7205 3145 7239 3179
rect 7573 3145 7607 3179
rect 7849 3145 7883 3179
rect 10793 3145 10827 3179
rect 11437 3145 11471 3179
rect 11805 3145 11839 3179
rect 12633 3145 12667 3179
rect 13093 3145 13127 3179
rect 1961 3077 1995 3111
rect 4997 3077 5031 3111
rect 4077 3009 4111 3043
rect 5549 3077 5583 3111
rect 6653 3009 6687 3043
rect 9321 3077 9355 3111
rect 9413 3009 9447 3043
rect 1777 2941 1811 2975
rect 4353 2941 4387 2975
rect 4815 2941 4849 2975
rect 5181 2941 5215 2975
rect 5365 2941 5399 2975
rect 5733 2941 5767 2975
rect 5917 2941 5951 2975
rect 6745 2941 6779 2975
rect 7083 2941 7117 2975
rect 7481 2941 7515 2975
rect 7573 2941 7607 2975
rect 8217 2941 8251 2975
rect 8401 2941 8435 2975
rect 8861 2941 8895 2975
rect 9045 2941 9079 2975
rect 9764 2941 9798 2975
rect 9960 2941 9994 2975
rect 10149 2941 10183 2975
rect 10333 2941 10367 2975
rect 11069 2941 11103 2975
rect 11161 2941 11195 2975
rect 11437 2941 11471 2975
rect 11937 2941 11971 2975
rect 12357 2941 12391 2975
rect 12817 2941 12851 2975
rect 13277 2941 13311 2975
rect 1593 2873 1627 2907
rect 3801 2873 3835 2907
rect 7757 2873 7791 2907
rect 8585 2873 8619 2907
rect 10057 2873 10091 2907
rect 11345 2873 11379 2907
rect 12081 2873 12115 2907
rect 12173 2873 12207 2907
rect 2329 2805 2363 2839
rect 4813 2805 4847 2839
rect 10977 2805 11011 2839
rect 2053 2601 2087 2635
rect 5365 2601 5399 2635
rect 5549 2601 5583 2635
rect 7113 2601 7147 2635
rect 10517 2601 10551 2635
rect 13093 2601 13127 2635
rect 3065 2533 3099 2567
rect 3525 2533 3559 2567
rect 4261 2533 4295 2567
rect 5273 2533 5307 2567
rect 7941 2533 7975 2567
rect 9873 2533 9907 2567
rect 1869 2465 1903 2499
rect 2329 2465 2363 2499
rect 2513 2465 2547 2499
rect 3249 2465 3283 2499
rect 3433 2465 3467 2499
rect 4164 2465 4198 2499
rect 4353 2465 4387 2499
rect 4537 2465 4571 2499
rect 5181 2465 5215 2499
rect 6193 2465 6227 2499
rect 6469 2465 6503 2499
rect 6617 2465 6651 2499
rect 6745 2465 6779 2499
rect 7021 2465 7055 2499
rect 7752 2465 7786 2499
rect 7849 2465 7883 2499
rect 8125 2465 8159 2499
rect 8493 2465 8527 2499
rect 8677 2465 8711 2499
rect 9505 2465 9539 2499
rect 10149 2465 10183 2499
rect 2697 2397 2731 2431
rect 6377 2397 6411 2431
rect 6837 2397 6871 2431
rect 9321 2397 9355 2431
rect 10057 2397 10091 2431
rect 3985 2329 4019 2363
rect 4997 2329 5031 2363
rect 10977 2533 11011 2567
rect 10609 2465 10643 2499
rect 10793 2465 10827 2499
rect 11345 2465 11379 2499
rect 11621 2397 11655 2431
rect 8677 2329 8711 2363
rect 10517 2329 10551 2363
rect 6009 2261 6043 2295
rect 6377 2261 6411 2295
rect 7573 2261 7607 2295
rect 2145 2057 2179 2091
rect 6653 2057 6687 2091
rect 7113 2057 7147 2091
rect 9229 2057 9263 2091
rect 9873 2057 9907 2091
rect 11253 2057 11287 2091
rect 13185 2057 13219 2091
rect 10425 1989 10459 2023
rect 11529 1989 11563 2023
rect 12265 1989 12299 2023
rect 3893 1921 3927 1955
rect 4813 1921 4847 1955
rect 8585 1921 8619 1955
rect 8861 1921 8895 1955
rect 9045 1921 9079 1955
rect 4537 1853 4571 1887
rect 4721 1853 4755 1887
rect 4906 1853 4940 1887
rect 5089 1853 5123 1887
rect 5641 1853 5675 1887
rect 5917 1853 5951 1887
rect 6101 1853 6135 1887
rect 6745 1853 6779 1887
rect 3617 1785 3651 1819
rect 4353 1785 4387 1819
rect 5733 1785 5767 1819
rect 5825 1785 5859 1819
rect 9137 1853 9171 1887
rect 10055 1853 10089 1887
rect 10517 1853 10551 1887
rect 11161 1853 11195 1887
rect 11529 1853 11563 1887
rect 11713 1853 11747 1887
rect 11989 1853 12023 1887
rect 12086 1853 12120 1887
rect 12817 1853 12851 1887
rect 13093 1853 13127 1887
rect 10977 1785 11011 1819
rect 11897 1785 11931 1819
rect 5457 1717 5491 1751
rect 9045 1717 9079 1751
rect 10057 1717 10091 1751
rect 12633 1717 12667 1751
rect 2421 1513 2455 1547
rect 2881 1513 2915 1547
rect 6101 1513 6135 1547
rect 6653 1513 6687 1547
rect 8769 1513 8803 1547
rect 9229 1513 9263 1547
rect 9781 1513 9815 1547
rect 11713 1513 11747 1547
rect 11897 1513 11931 1547
rect 12541 1513 12575 1547
rect 7297 1445 7331 1479
rect 2237 1377 2271 1411
rect 2697 1377 2731 1411
rect 3341 1377 3375 1411
rect 3525 1377 3559 1411
rect 3985 1377 4019 1411
rect 4077 1377 4111 1411
rect 6745 1377 6779 1411
rect 9413 1377 9447 1411
rect 11529 1377 11563 1411
rect 11713 1377 11747 1411
rect 12081 1377 12115 1411
rect 12357 1377 12391 1411
rect 4353 1309 4387 1343
rect 4629 1309 4663 1343
rect 7021 1309 7055 1343
rect 11253 1309 11287 1343
rect 3433 1241 3467 1275
<< metal1 >>
rect 1104 15802 13892 15824
rect 1104 15750 8246 15802
rect 8298 15750 8310 15802
rect 8362 15750 8374 15802
rect 8426 15750 8438 15802
rect 8490 15750 13892 15802
rect 1104 15728 13892 15750
rect 4614 15648 4620 15700
rect 4672 15688 4678 15700
rect 4893 15691 4951 15697
rect 4893 15688 4905 15691
rect 4672 15660 4905 15688
rect 4672 15648 4678 15660
rect 4893 15657 4905 15660
rect 4939 15657 4951 15691
rect 4893 15651 4951 15657
rect 4801 15623 4859 15629
rect 4801 15589 4813 15623
rect 4847 15620 4859 15623
rect 4982 15620 4988 15632
rect 4847 15592 4988 15620
rect 4847 15589 4859 15592
rect 4801 15583 4859 15589
rect 4982 15580 4988 15592
rect 5040 15580 5046 15632
rect 4157 15555 4215 15561
rect 4157 15521 4169 15555
rect 4203 15552 4215 15555
rect 4203 15524 4844 15552
rect 4203 15521 4215 15524
rect 4157 15515 4215 15521
rect 4816 15496 4844 15524
rect 4890 15512 4896 15564
rect 4948 15552 4954 15564
rect 5629 15555 5687 15561
rect 5629 15552 5641 15555
rect 4948 15524 5641 15552
rect 4948 15512 4954 15524
rect 5629 15521 5641 15524
rect 5675 15521 5687 15555
rect 5629 15515 5687 15521
rect 6181 15555 6239 15561
rect 6181 15521 6193 15555
rect 6227 15552 6239 15555
rect 6546 15552 6552 15564
rect 6227 15524 6552 15552
rect 6227 15521 6239 15524
rect 6181 15515 6239 15521
rect 6546 15512 6552 15524
rect 6604 15512 6610 15564
rect 6822 15552 6828 15564
rect 6783 15524 6828 15552
rect 6822 15512 6828 15524
rect 6880 15512 6886 15564
rect 7469 15555 7527 15561
rect 7469 15521 7481 15555
rect 7515 15521 7527 15555
rect 7469 15515 7527 15521
rect 4798 15444 4804 15496
rect 4856 15444 4862 15496
rect 5077 15487 5135 15493
rect 5077 15453 5089 15487
rect 5123 15484 5135 15487
rect 5810 15484 5816 15496
rect 5123 15456 5816 15484
rect 5123 15453 5135 15456
rect 5077 15447 5135 15453
rect 5810 15444 5816 15456
rect 5868 15444 5874 15496
rect 6454 15444 6460 15496
rect 6512 15484 6518 15496
rect 7484 15484 7512 15515
rect 8754 15512 8760 15564
rect 8812 15552 8818 15564
rect 9401 15555 9459 15561
rect 9401 15552 9413 15555
rect 8812 15524 9413 15552
rect 8812 15512 8818 15524
rect 9401 15521 9413 15524
rect 9447 15521 9459 15555
rect 10226 15552 10232 15564
rect 10187 15524 10232 15552
rect 9401 15515 9459 15521
rect 10226 15512 10232 15524
rect 10284 15512 10290 15564
rect 8018 15484 8024 15496
rect 6512 15456 7512 15484
rect 7979 15456 8024 15484
rect 6512 15444 6518 15456
rect 8018 15444 8024 15456
rect 8076 15444 8082 15496
rect 8573 15487 8631 15493
rect 8573 15453 8585 15487
rect 8619 15453 8631 15487
rect 8573 15447 8631 15453
rect 6089 15419 6147 15425
rect 6089 15385 6101 15419
rect 6135 15416 6147 15419
rect 7006 15416 7012 15428
rect 6135 15388 7012 15416
rect 6135 15385 6147 15388
rect 6089 15379 6147 15385
rect 7006 15376 7012 15388
rect 7064 15376 7070 15428
rect 8481 15419 8539 15425
rect 8481 15385 8493 15419
rect 8527 15385 8539 15419
rect 8588 15416 8616 15447
rect 9217 15419 9275 15425
rect 9217 15416 9229 15419
rect 8588 15388 9229 15416
rect 8481 15379 8539 15385
rect 9217 15385 9229 15388
rect 9263 15385 9275 15419
rect 9217 15379 9275 15385
rect 4062 15348 4068 15360
rect 4023 15320 4068 15348
rect 4062 15308 4068 15320
rect 4120 15308 4126 15360
rect 4433 15351 4491 15357
rect 4433 15317 4445 15351
rect 4479 15348 4491 15351
rect 4614 15348 4620 15360
rect 4479 15320 4620 15348
rect 4479 15317 4491 15320
rect 4433 15311 4491 15317
rect 4614 15308 4620 15320
rect 4672 15308 4678 15360
rect 5442 15348 5448 15360
rect 5403 15320 5448 15348
rect 5442 15308 5448 15320
rect 5500 15308 5506 15360
rect 6638 15348 6644 15360
rect 6599 15320 6644 15348
rect 6638 15308 6644 15320
rect 6696 15308 6702 15360
rect 7282 15348 7288 15360
rect 7243 15320 7288 15348
rect 7282 15308 7288 15320
rect 7340 15308 7346 15360
rect 8496 15348 8524 15379
rect 8570 15348 8576 15360
rect 8496 15320 8576 15348
rect 8570 15308 8576 15320
rect 8628 15308 8634 15360
rect 10134 15348 10140 15360
rect 10095 15320 10140 15348
rect 10134 15308 10140 15320
rect 10192 15308 10198 15360
rect 1104 15258 13892 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 12246 15258
rect 12298 15206 12310 15258
rect 12362 15206 12374 15258
rect 12426 15206 12438 15258
rect 12490 15206 13892 15258
rect 1104 15184 13892 15206
rect 5994 15144 6000 15156
rect 5955 15116 6000 15144
rect 5994 15104 6000 15116
rect 6052 15104 6058 15156
rect 10410 15144 10416 15156
rect 10152 15116 10416 15144
rect 6914 14968 6920 15020
rect 6972 15008 6978 15020
rect 7193 15011 7251 15017
rect 7193 15008 7205 15011
rect 6972 14980 7205 15008
rect 6972 14968 6978 14980
rect 7193 14977 7205 14980
rect 7239 14977 7251 15011
rect 7193 14971 7251 14977
rect 7377 15011 7435 15017
rect 7377 14977 7389 15011
rect 7423 15008 7435 15011
rect 7926 15008 7932 15020
rect 7423 14980 7932 15008
rect 7423 14977 7435 14980
rect 7377 14971 7435 14977
rect 7926 14968 7932 14980
rect 7984 15008 7990 15020
rect 8478 15008 8484 15020
rect 7984 14980 8484 15008
rect 7984 14968 7990 14980
rect 8478 14968 8484 14980
rect 8536 14968 8542 15020
rect 9858 15008 9864 15020
rect 9819 14980 9864 15008
rect 9858 14968 9864 14980
rect 9916 14968 9922 15020
rect 10045 15011 10103 15017
rect 10045 14977 10057 15011
rect 10091 15008 10103 15011
rect 10152 15008 10180 15116
rect 10410 15104 10416 15116
rect 10468 15144 10474 15156
rect 10468 15116 10732 15144
rect 10468 15104 10474 15116
rect 10597 15079 10655 15085
rect 10597 15045 10609 15079
rect 10643 15045 10655 15079
rect 10597 15039 10655 15045
rect 10091 14980 10180 15008
rect 10091 14977 10103 14980
rect 10045 14971 10103 14977
rect 3789 14943 3847 14949
rect 3789 14909 3801 14943
rect 3835 14940 3847 14943
rect 4614 14940 4620 14952
rect 3835 14912 4620 14940
rect 3835 14909 3847 14912
rect 3789 14903 3847 14909
rect 4614 14900 4620 14912
rect 4672 14900 4678 14952
rect 4709 14943 4767 14949
rect 4709 14909 4721 14943
rect 4755 14940 4767 14943
rect 4890 14940 4896 14952
rect 4755 14912 4896 14940
rect 4755 14909 4767 14912
rect 4709 14903 4767 14909
rect 4890 14900 4896 14912
rect 4948 14900 4954 14952
rect 5997 14943 6055 14949
rect 5997 14909 6009 14943
rect 6043 14940 6055 14943
rect 6638 14940 6644 14952
rect 6043 14912 6644 14940
rect 6043 14909 6055 14912
rect 5997 14903 6055 14909
rect 6638 14900 6644 14912
rect 6696 14900 6702 14952
rect 7837 14943 7895 14949
rect 7837 14909 7849 14943
rect 7883 14940 7895 14943
rect 8018 14940 8024 14952
rect 7883 14912 8024 14940
rect 7883 14909 7895 14912
rect 7837 14903 7895 14909
rect 8018 14900 8024 14912
rect 8076 14940 8082 14952
rect 10612 14940 10640 15039
rect 10704 15008 10732 15116
rect 11149 15011 11207 15017
rect 11149 15008 11161 15011
rect 10704 14980 11161 15008
rect 11149 14977 11161 14980
rect 11195 14977 11207 15011
rect 11149 14971 11207 14977
rect 8076 14912 10640 14940
rect 11057 14943 11115 14949
rect 8076 14900 8082 14912
rect 11057 14909 11069 14943
rect 11103 14940 11115 14943
rect 12526 14940 12532 14952
rect 11103 14912 12532 14940
rect 11103 14909 11115 14912
rect 11057 14903 11115 14909
rect 12526 14900 12532 14912
rect 12584 14900 12590 14952
rect 4525 14875 4583 14881
rect 4525 14841 4537 14875
rect 4571 14841 4583 14875
rect 8570 14872 8576 14884
rect 8531 14844 8576 14872
rect 4525 14835 4583 14841
rect 4540 14804 4568 14835
rect 8570 14832 8576 14844
rect 8628 14832 8634 14884
rect 8754 14872 8760 14884
rect 8715 14844 8760 14872
rect 8754 14832 8760 14844
rect 8812 14832 8818 14884
rect 4798 14804 4804 14816
rect 4540 14776 4804 14804
rect 4798 14764 4804 14776
rect 4856 14764 4862 14816
rect 6730 14804 6736 14816
rect 6691 14776 6736 14804
rect 6730 14764 6736 14776
rect 6788 14764 6794 14816
rect 7101 14807 7159 14813
rect 7101 14773 7113 14807
rect 7147 14804 7159 14807
rect 8018 14804 8024 14816
rect 7147 14776 8024 14804
rect 7147 14773 7159 14776
rect 7101 14767 7159 14773
rect 8018 14764 8024 14776
rect 8076 14764 8082 14816
rect 9214 14764 9220 14816
rect 9272 14804 9278 14816
rect 9401 14807 9459 14813
rect 9401 14804 9413 14807
rect 9272 14776 9413 14804
rect 9272 14764 9278 14776
rect 9401 14773 9413 14776
rect 9447 14773 9459 14807
rect 9766 14804 9772 14816
rect 9727 14776 9772 14804
rect 9401 14767 9459 14773
rect 9766 14764 9772 14776
rect 9824 14764 9830 14816
rect 10965 14807 11023 14813
rect 10965 14773 10977 14807
rect 11011 14804 11023 14807
rect 11146 14804 11152 14816
rect 11011 14776 11152 14804
rect 11011 14773 11023 14776
rect 10965 14767 11023 14773
rect 11146 14764 11152 14776
rect 11204 14764 11210 14816
rect 1104 14714 13892 14736
rect 1104 14662 8246 14714
rect 8298 14662 8310 14714
rect 8362 14662 8374 14714
rect 8426 14662 8438 14714
rect 8490 14662 13892 14714
rect 1104 14640 13892 14662
rect 1854 14560 1860 14612
rect 1912 14600 1918 14612
rect 2225 14603 2283 14609
rect 2225 14600 2237 14603
rect 1912 14572 2237 14600
rect 1912 14560 1918 14572
rect 2225 14569 2237 14572
rect 2271 14569 2283 14603
rect 2225 14563 2283 14569
rect 8570 14560 8576 14612
rect 8628 14600 8634 14612
rect 11057 14603 11115 14609
rect 11057 14600 11069 14603
rect 8628 14572 11069 14600
rect 8628 14560 8634 14572
rect 11057 14569 11069 14572
rect 11103 14569 11115 14603
rect 11057 14563 11115 14569
rect 3881 14535 3939 14541
rect 3881 14501 3893 14535
rect 3927 14532 3939 14535
rect 4062 14532 4068 14544
rect 3927 14504 4068 14532
rect 3927 14501 3939 14504
rect 3881 14495 3939 14501
rect 4062 14492 4068 14504
rect 4120 14492 4126 14544
rect 4798 14492 4804 14544
rect 4856 14532 4862 14544
rect 5169 14535 5227 14541
rect 5169 14532 5181 14535
rect 4856 14504 5181 14532
rect 4856 14492 4862 14504
rect 5169 14501 5181 14504
rect 5215 14501 5227 14535
rect 5169 14495 5227 14501
rect 5261 14535 5319 14541
rect 5261 14501 5273 14535
rect 5307 14532 5319 14535
rect 5442 14532 5448 14544
rect 5307 14504 5448 14532
rect 5307 14501 5319 14504
rect 5261 14495 5319 14501
rect 5442 14492 5448 14504
rect 5500 14492 5506 14544
rect 7282 14492 7288 14544
rect 7340 14532 7346 14544
rect 7377 14535 7435 14541
rect 7377 14532 7389 14535
rect 7340 14504 7389 14532
rect 7340 14492 7346 14504
rect 7377 14501 7389 14504
rect 7423 14501 7435 14535
rect 7377 14495 7435 14501
rect 2133 14467 2191 14473
rect 2133 14433 2145 14467
rect 2179 14464 2191 14467
rect 3050 14464 3056 14476
rect 2179 14436 3056 14464
rect 2179 14433 2191 14436
rect 2133 14427 2191 14433
rect 3050 14424 3056 14436
rect 3108 14424 3114 14476
rect 3145 14467 3203 14473
rect 3145 14433 3157 14467
rect 3191 14433 3203 14467
rect 3145 14427 3203 14433
rect 2038 14356 2044 14408
rect 2096 14396 2102 14408
rect 2317 14399 2375 14405
rect 2317 14396 2329 14399
rect 2096 14368 2329 14396
rect 2096 14356 2102 14368
rect 2317 14365 2329 14368
rect 2363 14365 2375 14399
rect 2317 14359 2375 14365
rect 2774 14288 2780 14340
rect 2832 14328 2838 14340
rect 2961 14331 3019 14337
rect 2961 14328 2973 14331
rect 2832 14300 2973 14328
rect 2832 14288 2838 14300
rect 2961 14297 2973 14300
rect 3007 14297 3019 14331
rect 2961 14291 3019 14297
rect 1762 14260 1768 14272
rect 1723 14232 1768 14260
rect 1762 14220 1768 14232
rect 1820 14220 1826 14272
rect 3160 14260 3188 14427
rect 4614 14424 4620 14476
rect 4672 14464 4678 14476
rect 4709 14467 4767 14473
rect 4709 14464 4721 14467
rect 4672 14436 4721 14464
rect 4672 14424 4678 14436
rect 4709 14433 4721 14436
rect 4755 14433 4767 14467
rect 4709 14427 4767 14433
rect 5537 14467 5595 14473
rect 5537 14433 5549 14467
rect 5583 14464 5595 14467
rect 5902 14464 5908 14476
rect 5583 14436 5908 14464
rect 5583 14433 5595 14436
rect 5537 14427 5595 14433
rect 5902 14424 5908 14436
rect 5960 14424 5966 14476
rect 6454 14464 6460 14476
rect 6415 14436 6460 14464
rect 6454 14424 6460 14436
rect 6512 14424 6518 14476
rect 6546 14424 6552 14476
rect 6604 14464 6610 14476
rect 7469 14467 7527 14473
rect 7469 14464 7481 14467
rect 6604 14436 7481 14464
rect 6604 14424 6610 14436
rect 7469 14433 7481 14436
rect 7515 14433 7527 14467
rect 7469 14427 7527 14433
rect 7558 14424 7564 14476
rect 7616 14464 7622 14476
rect 8205 14467 8263 14473
rect 8205 14464 8217 14467
rect 7616 14436 8217 14464
rect 7616 14424 7622 14436
rect 8205 14433 8217 14436
rect 8251 14433 8263 14467
rect 8846 14464 8852 14476
rect 8205 14427 8263 14433
rect 8312 14436 8852 14464
rect 3326 14356 3332 14408
rect 3384 14396 3390 14408
rect 4433 14399 4491 14405
rect 4433 14396 4445 14399
rect 3384 14368 4445 14396
rect 3384 14356 3390 14368
rect 4433 14365 4445 14368
rect 4479 14396 4491 14399
rect 6730 14396 6736 14408
rect 4479 14368 6736 14396
rect 4479 14365 4491 14368
rect 4433 14359 4491 14365
rect 6730 14356 6736 14368
rect 6788 14356 6794 14408
rect 7929 14399 7987 14405
rect 7929 14365 7941 14399
rect 7975 14396 7987 14399
rect 8312 14396 8340 14436
rect 8846 14424 8852 14436
rect 8904 14424 8910 14476
rect 9214 14464 9220 14476
rect 9175 14436 9220 14464
rect 9214 14424 9220 14436
rect 9272 14424 9278 14476
rect 10689 14467 10747 14473
rect 10689 14433 10701 14467
rect 10735 14464 10747 14467
rect 10962 14464 10968 14476
rect 10735 14436 10968 14464
rect 10735 14433 10747 14436
rect 10689 14427 10747 14433
rect 10962 14424 10968 14436
rect 11020 14464 11026 14476
rect 11701 14467 11759 14473
rect 11701 14464 11713 14467
rect 11020 14436 11713 14464
rect 11020 14424 11026 14436
rect 11701 14433 11713 14436
rect 11747 14433 11759 14467
rect 11701 14427 11759 14433
rect 7975 14368 8340 14396
rect 8757 14399 8815 14405
rect 7975 14365 7987 14368
rect 7929 14359 7987 14365
rect 8757 14365 8769 14399
rect 8803 14396 8815 14399
rect 11149 14399 11207 14405
rect 11149 14396 11161 14399
rect 8803 14368 11161 14396
rect 8803 14365 8815 14368
rect 8757 14359 8815 14365
rect 11149 14365 11161 14368
rect 11195 14365 11207 14399
rect 11149 14359 11207 14365
rect 3878 14288 3884 14340
rect 3936 14328 3942 14340
rect 3973 14331 4031 14337
rect 3973 14328 3985 14331
rect 3936 14300 3985 14328
rect 3936 14288 3942 14300
rect 3973 14297 3985 14300
rect 4019 14297 4031 14331
rect 6822 14328 6828 14340
rect 6783 14300 6828 14328
rect 3973 14291 4031 14297
rect 6822 14288 6828 14300
rect 6880 14288 6886 14340
rect 8662 14328 8668 14340
rect 8623 14300 8668 14328
rect 8662 14288 8668 14300
rect 8720 14288 8726 14340
rect 10505 14331 10563 14337
rect 10505 14297 10517 14331
rect 10551 14297 10563 14331
rect 10505 14291 10563 14297
rect 9950 14260 9956 14272
rect 3160 14232 9956 14260
rect 9950 14220 9956 14232
rect 10008 14260 10014 14272
rect 10520 14260 10548 14291
rect 10008 14232 10548 14260
rect 10008 14220 10014 14232
rect 10870 14220 10876 14272
rect 10928 14260 10934 14272
rect 11517 14263 11575 14269
rect 11517 14260 11529 14263
rect 10928 14232 11529 14260
rect 10928 14220 10934 14232
rect 11517 14229 11529 14232
rect 11563 14229 11575 14263
rect 11517 14223 11575 14229
rect 1104 14170 13892 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 12246 14170
rect 12298 14118 12310 14170
rect 12362 14118 12374 14170
rect 12426 14118 12438 14170
rect 12490 14118 13892 14170
rect 1104 14096 13892 14118
rect 5902 14056 5908 14068
rect 5863 14028 5908 14056
rect 5902 14016 5908 14028
rect 5960 14016 5966 14068
rect 8662 14016 8668 14068
rect 8720 14056 8726 14068
rect 8720 14028 12434 14056
rect 8720 14016 8726 14028
rect 4062 13948 4068 14000
rect 4120 13988 4126 14000
rect 4120 13960 5488 13988
rect 4120 13948 4126 13960
rect 3878 13880 3884 13932
rect 3936 13920 3942 13932
rect 5460 13929 5488 13960
rect 4893 13923 4951 13929
rect 4893 13920 4905 13923
rect 3936 13892 4905 13920
rect 3936 13880 3942 13892
rect 4893 13889 4905 13892
rect 4939 13889 4951 13923
rect 4893 13883 4951 13889
rect 5353 13923 5411 13929
rect 5353 13889 5365 13923
rect 5399 13889 5411 13923
rect 5353 13883 5411 13889
rect 5445 13923 5503 13929
rect 5445 13889 5457 13923
rect 5491 13889 5503 13923
rect 5920 13920 5948 14016
rect 6822 13948 6828 14000
rect 6880 13988 6886 14000
rect 6917 13991 6975 13997
rect 6917 13988 6929 13991
rect 6880 13960 6929 13988
rect 6880 13948 6886 13960
rect 6917 13957 6929 13960
rect 6963 13988 6975 13991
rect 8570 13988 8576 14000
rect 6963 13960 8576 13988
rect 6963 13957 6975 13960
rect 6917 13951 6975 13957
rect 8570 13948 8576 13960
rect 8628 13948 8634 14000
rect 9048 13997 9076 14028
rect 9033 13991 9091 13997
rect 9033 13957 9045 13991
rect 9079 13957 9091 13991
rect 9950 13988 9956 14000
rect 9911 13960 9956 13988
rect 9033 13951 9091 13957
rect 9950 13948 9956 13960
rect 10008 13948 10014 14000
rect 10226 13948 10232 14000
rect 10284 13988 10290 14000
rect 10781 13991 10839 13997
rect 10781 13988 10793 13991
rect 10284 13960 10793 13988
rect 10284 13948 10290 13960
rect 10781 13957 10793 13960
rect 10827 13957 10839 13991
rect 10781 13951 10839 13957
rect 11698 13948 11704 14000
rect 11756 13988 11762 14000
rect 12253 13991 12311 13997
rect 12253 13988 12265 13991
rect 11756 13960 12265 13988
rect 11756 13948 11762 13960
rect 12253 13957 12265 13960
rect 12299 13957 12311 13991
rect 12253 13951 12311 13957
rect 6457 13923 6515 13929
rect 6457 13920 6469 13923
rect 5920 13892 6469 13920
rect 5445 13883 5503 13889
rect 6457 13889 6469 13892
rect 6503 13889 6515 13923
rect 7006 13920 7012 13932
rect 6967 13892 7012 13920
rect 6457 13883 6515 13889
rect 1762 13812 1768 13864
rect 1820 13852 1826 13864
rect 1857 13855 1915 13861
rect 1857 13852 1869 13855
rect 1820 13824 1869 13852
rect 1820 13812 1826 13824
rect 1857 13821 1869 13824
rect 1903 13821 1915 13855
rect 3326 13852 3332 13864
rect 3287 13824 3332 13852
rect 1857 13815 1915 13821
rect 3326 13812 3332 13824
rect 3384 13812 3390 13864
rect 4798 13852 4804 13864
rect 4759 13824 4804 13852
rect 4798 13812 4804 13824
rect 4856 13812 4862 13864
rect 5368 13852 5396 13883
rect 7006 13880 7012 13892
rect 7064 13880 7070 13932
rect 9214 13880 9220 13932
rect 9272 13920 9278 13932
rect 9493 13923 9551 13929
rect 9493 13920 9505 13923
rect 9272 13892 9505 13920
rect 9272 13880 9278 13892
rect 9493 13889 9505 13892
rect 9539 13889 9551 13923
rect 9493 13883 9551 13889
rect 10045 13923 10103 13929
rect 10045 13889 10057 13923
rect 10091 13920 10103 13923
rect 10134 13920 10140 13932
rect 10091 13892 10140 13920
rect 10091 13889 10103 13892
rect 10045 13883 10103 13889
rect 10134 13880 10140 13892
rect 10192 13880 10198 13932
rect 10870 13920 10876 13932
rect 10831 13892 10876 13920
rect 10870 13880 10876 13892
rect 10928 13880 10934 13932
rect 12406 13920 12434 14028
rect 12710 13920 12716 13932
rect 12406 13892 12716 13920
rect 12710 13880 12716 13892
rect 12768 13880 12774 13932
rect 5810 13852 5816 13864
rect 5368 13824 5816 13852
rect 5810 13812 5816 13824
rect 5868 13812 5874 13864
rect 7558 13852 7564 13864
rect 7519 13824 7564 13852
rect 7558 13812 7564 13824
rect 7616 13812 7622 13864
rect 8754 13852 8760 13864
rect 8715 13824 8760 13852
rect 8754 13812 8760 13824
rect 8812 13812 8818 13864
rect 10318 13852 10324 13864
rect 10279 13824 10324 13852
rect 10318 13812 10324 13824
rect 10376 13812 10382 13864
rect 10962 13812 10968 13864
rect 11020 13852 11026 13864
rect 11701 13855 11759 13861
rect 11701 13852 11713 13855
rect 11020 13824 11713 13852
rect 11020 13812 11026 13824
rect 11701 13821 11713 13824
rect 11747 13821 11759 13855
rect 12434 13852 12440 13864
rect 12395 13824 12440 13852
rect 11701 13815 11759 13821
rect 12434 13812 12440 13824
rect 12492 13812 12498 13864
rect 13173 13855 13231 13861
rect 13173 13821 13185 13855
rect 13219 13852 13231 13855
rect 13262 13852 13268 13864
rect 13219 13824 13268 13852
rect 13219 13821 13231 13824
rect 13173 13815 13231 13821
rect 13262 13812 13268 13824
rect 13320 13812 13326 13864
rect 2498 13784 2504 13796
rect 2459 13756 2504 13784
rect 2498 13744 2504 13756
rect 2556 13744 2562 13796
rect 2774 13744 2780 13796
rect 2832 13784 2838 13796
rect 11882 13784 11888 13796
rect 2832 13756 2877 13784
rect 11843 13756 11888 13784
rect 2832 13744 2838 13756
rect 11882 13744 11888 13756
rect 11940 13744 11946 13796
rect 5534 13716 5540 13728
rect 5495 13688 5540 13716
rect 5534 13676 5540 13688
rect 5592 13676 5598 13728
rect 11238 13716 11244 13728
rect 11199 13688 11244 13716
rect 11238 13676 11244 13688
rect 11296 13676 11302 13728
rect 11333 13719 11391 13725
rect 11333 13685 11345 13719
rect 11379 13716 11391 13719
rect 11606 13716 11612 13728
rect 11379 13688 11612 13716
rect 11379 13685 11391 13688
rect 11333 13679 11391 13685
rect 11606 13676 11612 13688
rect 11664 13676 11670 13728
rect 12986 13716 12992 13728
rect 12947 13688 12992 13716
rect 12986 13676 12992 13688
rect 13044 13676 13050 13728
rect 1104 13626 13892 13648
rect 1104 13574 8246 13626
rect 8298 13574 8310 13626
rect 8362 13574 8374 13626
rect 8426 13574 8438 13626
rect 8490 13574 13892 13626
rect 1104 13552 13892 13574
rect 2866 13512 2872 13524
rect 2827 13484 2872 13512
rect 2866 13472 2872 13484
rect 2924 13472 2930 13524
rect 3050 13472 3056 13524
rect 3108 13512 3114 13524
rect 3881 13515 3939 13521
rect 3881 13512 3893 13515
rect 3108 13484 3893 13512
rect 3108 13472 3114 13484
rect 3881 13481 3893 13484
rect 3927 13481 3939 13515
rect 8846 13512 8852 13524
rect 3881 13475 3939 13481
rect 7576 13484 8852 13512
rect 1673 13447 1731 13453
rect 1673 13413 1685 13447
rect 1719 13444 1731 13447
rect 2409 13447 2467 13453
rect 2409 13444 2421 13447
rect 1719 13416 2421 13444
rect 1719 13413 1731 13416
rect 1673 13407 1731 13413
rect 2409 13413 2421 13416
rect 2455 13444 2467 13447
rect 2498 13444 2504 13456
rect 2455 13416 2504 13444
rect 2455 13413 2467 13416
rect 2409 13407 2467 13413
rect 2498 13404 2504 13416
rect 2556 13404 2562 13456
rect 4617 13447 4675 13453
rect 4617 13413 4629 13447
rect 4663 13444 4675 13447
rect 4798 13444 4804 13456
rect 4663 13416 4804 13444
rect 4663 13413 4675 13416
rect 4617 13407 4675 13413
rect 4798 13404 4804 13416
rect 4856 13404 4862 13456
rect 5169 13447 5227 13453
rect 5169 13413 5181 13447
rect 5215 13444 5227 13447
rect 6362 13444 6368 13456
rect 5215 13416 6368 13444
rect 5215 13413 5227 13416
rect 5169 13407 5227 13413
rect 6362 13404 6368 13416
rect 6420 13404 6426 13456
rect 6546 13404 6552 13456
rect 6604 13444 6610 13456
rect 6825 13447 6883 13453
rect 6825 13444 6837 13447
rect 6604 13416 6837 13444
rect 6604 13404 6610 13416
rect 6825 13413 6837 13416
rect 6871 13413 6883 13447
rect 6825 13407 6883 13413
rect 1762 13336 1768 13388
rect 1820 13376 1826 13388
rect 1949 13379 2007 13385
rect 1949 13376 1961 13379
rect 1820 13348 1961 13376
rect 1820 13336 1826 13348
rect 1949 13345 1961 13348
rect 1995 13345 2007 13379
rect 1949 13339 2007 13345
rect 2961 13379 3019 13385
rect 2961 13345 2973 13379
rect 3007 13376 3019 13379
rect 3050 13376 3056 13388
rect 3007 13348 3056 13376
rect 3007 13345 3019 13348
rect 2961 13339 3019 13345
rect 3050 13336 3056 13348
rect 3108 13336 3114 13388
rect 3513 13379 3571 13385
rect 3513 13345 3525 13379
rect 3559 13345 3571 13379
rect 3513 13339 3571 13345
rect 4065 13379 4123 13385
rect 4065 13345 4077 13379
rect 4111 13345 4123 13379
rect 4065 13339 4123 13345
rect 4433 13379 4491 13385
rect 4433 13345 4445 13379
rect 4479 13376 4491 13379
rect 4706 13376 4712 13388
rect 4479 13348 4712 13376
rect 4479 13345 4491 13348
rect 4433 13339 4491 13345
rect 2501 13311 2559 13317
rect 2501 13277 2513 13311
rect 2547 13277 2559 13311
rect 2501 13271 2559 13277
rect 2516 13240 2544 13271
rect 2774 13268 2780 13320
rect 2832 13308 2838 13320
rect 3528 13308 3556 13339
rect 2832 13280 3556 13308
rect 4080 13308 4108 13339
rect 4706 13336 4712 13348
rect 4764 13336 4770 13388
rect 5350 13376 5356 13388
rect 5311 13348 5356 13376
rect 5350 13336 5356 13348
rect 5408 13336 5414 13388
rect 5718 13336 5724 13388
rect 5776 13376 5782 13388
rect 5813 13379 5871 13385
rect 5813 13376 5825 13379
rect 5776 13348 5825 13376
rect 5776 13336 5782 13348
rect 5813 13345 5825 13348
rect 5859 13345 5871 13379
rect 5813 13339 5871 13345
rect 5902 13336 5908 13388
rect 5960 13376 5966 13388
rect 5997 13379 6055 13385
rect 5997 13376 6009 13379
rect 5960 13348 6009 13376
rect 5960 13336 5966 13348
rect 5997 13345 6009 13348
rect 6043 13345 6055 13379
rect 5997 13339 6055 13345
rect 6454 13336 6460 13388
rect 6512 13376 6518 13388
rect 7576 13385 7604 13484
rect 8846 13472 8852 13484
rect 8904 13512 8910 13524
rect 9306 13512 9312 13524
rect 8904 13484 9312 13512
rect 8904 13472 8910 13484
rect 9306 13472 9312 13484
rect 9364 13472 9370 13524
rect 8481 13447 8539 13453
rect 8481 13413 8493 13447
rect 8527 13444 8539 13447
rect 8570 13444 8576 13456
rect 8527 13416 8576 13444
rect 8527 13413 8539 13416
rect 8481 13407 8539 13413
rect 8570 13404 8576 13416
rect 8628 13404 8634 13456
rect 8665 13447 8723 13453
rect 8665 13413 8677 13447
rect 8711 13444 8723 13447
rect 8754 13444 8760 13456
rect 8711 13416 8760 13444
rect 8711 13413 8723 13416
rect 8665 13407 8723 13413
rect 8754 13404 8760 13416
rect 8812 13404 8818 13456
rect 10226 13444 10232 13456
rect 10187 13416 10232 13444
rect 10226 13404 10232 13416
rect 10284 13404 10290 13456
rect 10505 13447 10563 13453
rect 10505 13413 10517 13447
rect 10551 13444 10563 13447
rect 10962 13444 10968 13456
rect 10551 13416 10968 13444
rect 10551 13413 10563 13416
rect 10505 13407 10563 13413
rect 10962 13404 10968 13416
rect 11020 13404 11026 13456
rect 11977 13447 12035 13453
rect 11977 13413 11989 13447
rect 12023 13444 12035 13447
rect 12434 13444 12440 13456
rect 12023 13416 12440 13444
rect 12023 13413 12035 13416
rect 11977 13407 12035 13413
rect 12434 13404 12440 13416
rect 12492 13444 12498 13456
rect 13170 13444 13176 13456
rect 12492 13416 13176 13444
rect 12492 13404 12498 13416
rect 13170 13404 13176 13416
rect 13228 13404 13234 13456
rect 6641 13379 6699 13385
rect 6641 13376 6653 13379
rect 6512 13348 6653 13376
rect 6512 13336 6518 13348
rect 6641 13345 6653 13348
rect 6687 13345 6699 13379
rect 6641 13339 6699 13345
rect 7561 13379 7619 13385
rect 7561 13345 7573 13379
rect 7607 13345 7619 13379
rect 7561 13339 7619 13345
rect 5166 13308 5172 13320
rect 4080 13280 5172 13308
rect 2832 13268 2838 13280
rect 5166 13268 5172 13280
rect 5224 13268 5230 13320
rect 6656 13308 6684 13339
rect 7650 13336 7656 13388
rect 7708 13376 7714 13388
rect 8021 13379 8079 13385
rect 8021 13376 8033 13379
rect 7708 13348 8033 13376
rect 7708 13336 7714 13348
rect 8021 13345 8033 13348
rect 8067 13345 8079 13379
rect 8021 13339 8079 13345
rect 8110 13336 8116 13388
rect 8168 13376 8174 13388
rect 9125 13379 9183 13385
rect 9125 13376 9137 13379
rect 8168 13348 9137 13376
rect 8168 13336 8174 13348
rect 9125 13345 9137 13348
rect 9171 13376 9183 13379
rect 9490 13376 9496 13388
rect 9171 13348 9496 13376
rect 9171 13345 9183 13348
rect 9125 13339 9183 13345
rect 9490 13336 9496 13348
rect 9548 13336 9554 13388
rect 9585 13379 9643 13385
rect 9585 13345 9597 13379
rect 9631 13376 9643 13379
rect 9674 13376 9680 13388
rect 9631 13348 9680 13376
rect 9631 13345 9643 13348
rect 9585 13339 9643 13345
rect 9674 13336 9680 13348
rect 9732 13376 9738 13388
rect 10318 13376 10324 13388
rect 9732 13348 10324 13376
rect 9732 13336 9738 13348
rect 10318 13336 10324 13348
rect 10376 13336 10382 13388
rect 11057 13379 11115 13385
rect 11057 13345 11069 13379
rect 11103 13345 11115 13379
rect 11057 13339 11115 13345
rect 7837 13311 7895 13317
rect 7837 13308 7849 13311
rect 6656 13280 7849 13308
rect 7837 13277 7849 13280
rect 7883 13277 7895 13311
rect 7837 13271 7895 13277
rect 7926 13268 7932 13320
rect 7984 13308 7990 13320
rect 8846 13308 8852 13320
rect 7984 13280 8852 13308
rect 7984 13268 7990 13280
rect 8846 13268 8852 13280
rect 8904 13308 8910 13320
rect 10410 13308 10416 13320
rect 8904 13280 10416 13308
rect 8904 13268 8910 13280
rect 10410 13268 10416 13280
rect 10468 13268 10474 13320
rect 3329 13243 3387 13249
rect 3329 13240 3341 13243
rect 2516 13212 3341 13240
rect 3329 13209 3341 13212
rect 3375 13209 3387 13243
rect 3329 13203 3387 13209
rect 7374 13200 7380 13252
rect 7432 13240 7438 13252
rect 11072 13240 11100 13339
rect 11606 13336 11612 13388
rect 11664 13376 11670 13388
rect 11701 13379 11759 13385
rect 11701 13376 11713 13379
rect 11664 13348 11713 13376
rect 11664 13336 11670 13348
rect 11701 13345 11713 13348
rect 11747 13345 11759 13379
rect 12710 13376 12716 13388
rect 12671 13348 12716 13376
rect 11701 13339 11759 13345
rect 12710 13336 12716 13348
rect 12768 13336 12774 13388
rect 12897 13379 12955 13385
rect 12897 13345 12909 13379
rect 12943 13376 12955 13379
rect 13354 13376 13360 13388
rect 12943 13348 13360 13376
rect 12943 13345 12955 13348
rect 12897 13339 12955 13345
rect 13354 13336 13360 13348
rect 13412 13336 13418 13388
rect 11330 13240 11336 13252
rect 7432 13212 11336 13240
rect 7432 13200 7438 13212
rect 11330 13200 11336 13212
rect 11388 13200 11394 13252
rect 1581 13175 1639 13181
rect 1581 13141 1593 13175
rect 1627 13172 1639 13175
rect 2958 13172 2964 13184
rect 1627 13144 2964 13172
rect 1627 13141 1639 13144
rect 1581 13135 1639 13141
rect 2958 13132 2964 13144
rect 3016 13132 3022 13184
rect 5074 13172 5080 13184
rect 5035 13144 5080 13172
rect 5074 13132 5080 13144
rect 5132 13132 5138 13184
rect 5721 13175 5779 13181
rect 5721 13141 5733 13175
rect 5767 13172 5779 13175
rect 6822 13172 6828 13184
rect 5767 13144 6828 13172
rect 5767 13141 5779 13144
rect 5721 13135 5779 13141
rect 6822 13132 6828 13144
rect 6880 13132 6886 13184
rect 9217 13175 9275 13181
rect 9217 13141 9229 13175
rect 9263 13172 9275 13175
rect 10962 13172 10968 13184
rect 9263 13144 10968 13172
rect 9263 13141 9275 13144
rect 9217 13135 9275 13141
rect 10962 13132 10968 13144
rect 11020 13132 11026 13184
rect 13078 13132 13084 13184
rect 13136 13172 13142 13184
rect 13173 13175 13231 13181
rect 13173 13172 13185 13175
rect 13136 13144 13185 13172
rect 13136 13132 13142 13144
rect 13173 13141 13185 13144
rect 13219 13141 13231 13175
rect 13173 13135 13231 13141
rect 1104 13082 13892 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 12246 13082
rect 12298 13030 12310 13082
rect 12362 13030 12374 13082
rect 12426 13030 12438 13082
rect 12490 13030 13892 13082
rect 1104 13008 13892 13030
rect 5074 12968 5080 12980
rect 2746 12940 5080 12968
rect 2038 12900 2044 12912
rect 1596 12872 2044 12900
rect 1596 12841 1624 12872
rect 2038 12860 2044 12872
rect 2096 12860 2102 12912
rect 1581 12835 1639 12841
rect 1581 12801 1593 12835
rect 1627 12801 1639 12835
rect 2746 12832 2774 12940
rect 5074 12928 5080 12940
rect 5132 12928 5138 12980
rect 5905 12971 5963 12977
rect 5905 12937 5917 12971
rect 5951 12968 5963 12971
rect 7558 12968 7564 12980
rect 5951 12940 7564 12968
rect 5951 12937 5963 12940
rect 5905 12931 5963 12937
rect 7558 12928 7564 12940
rect 7616 12928 7622 12980
rect 8018 12928 8024 12980
rect 8076 12968 8082 12980
rect 8205 12971 8263 12977
rect 8205 12968 8217 12971
rect 8076 12940 8217 12968
rect 8076 12928 8082 12940
rect 8205 12937 8217 12940
rect 8251 12968 8263 12971
rect 8938 12968 8944 12980
rect 8251 12940 8944 12968
rect 8251 12937 8263 12940
rect 8205 12931 8263 12937
rect 8938 12928 8944 12940
rect 8996 12928 9002 12980
rect 9674 12928 9680 12980
rect 9732 12968 9738 12980
rect 9769 12971 9827 12977
rect 9769 12968 9781 12971
rect 9732 12940 9781 12968
rect 9732 12928 9738 12940
rect 9769 12937 9781 12940
rect 9815 12937 9827 12971
rect 9769 12931 9827 12937
rect 2869 12903 2927 12909
rect 2869 12869 2881 12903
rect 2915 12900 2927 12903
rect 3050 12900 3056 12912
rect 2915 12872 3056 12900
rect 2915 12869 2927 12872
rect 2869 12863 2927 12869
rect 3050 12860 3056 12872
rect 3108 12860 3114 12912
rect 3234 12860 3240 12912
rect 3292 12900 3298 12912
rect 4338 12900 4344 12912
rect 3292 12872 4344 12900
rect 3292 12860 3298 12872
rect 4338 12860 4344 12872
rect 4396 12860 4402 12912
rect 6546 12860 6552 12912
rect 6604 12900 6610 12912
rect 9493 12903 9551 12909
rect 6604 12872 8984 12900
rect 6604 12860 6610 12872
rect 2958 12832 2964 12844
rect 1581 12795 1639 12801
rect 1780 12804 2774 12832
rect 2919 12804 2964 12832
rect 1780 12773 1808 12804
rect 2958 12792 2964 12804
rect 3016 12792 3022 12844
rect 3973 12835 4031 12841
rect 3973 12801 3985 12835
rect 4019 12832 4031 12835
rect 4706 12832 4712 12844
rect 4019 12804 4712 12832
rect 4019 12801 4031 12804
rect 3973 12795 4031 12801
rect 4706 12792 4712 12804
rect 4764 12792 4770 12844
rect 5353 12835 5411 12841
rect 5353 12801 5365 12835
rect 5399 12832 5411 12835
rect 5810 12832 5816 12844
rect 5399 12804 5816 12832
rect 5399 12801 5411 12804
rect 5353 12795 5411 12801
rect 5810 12792 5816 12804
rect 5868 12832 5874 12844
rect 6825 12835 6883 12841
rect 6825 12832 6837 12835
rect 5868 12804 6837 12832
rect 5868 12792 5874 12804
rect 6825 12801 6837 12804
rect 6871 12832 6883 12835
rect 8846 12832 8852 12844
rect 6871 12804 7420 12832
rect 8807 12804 8852 12832
rect 6871 12801 6883 12804
rect 6825 12795 6883 12801
rect 1765 12767 1823 12773
rect 1765 12733 1777 12767
rect 1811 12733 1823 12767
rect 2409 12767 2467 12773
rect 2409 12764 2421 12767
rect 1765 12727 1823 12733
rect 2148 12736 2421 12764
rect 2148 12640 2176 12736
rect 2409 12733 2421 12736
rect 2455 12733 2467 12767
rect 2409 12727 2467 12733
rect 3142 12724 3148 12776
rect 3200 12764 3206 12776
rect 3513 12767 3571 12773
rect 3513 12764 3525 12767
rect 3200 12736 3525 12764
rect 3200 12724 3206 12736
rect 3513 12733 3525 12736
rect 3559 12733 3571 12767
rect 3513 12727 3571 12733
rect 4525 12767 4583 12773
rect 4525 12733 4537 12767
rect 4571 12764 4583 12767
rect 5537 12767 5595 12773
rect 5537 12764 5549 12767
rect 4571 12736 5549 12764
rect 4571 12733 4583 12736
rect 4525 12727 4583 12733
rect 5537 12733 5549 12736
rect 5583 12733 5595 12767
rect 5537 12727 5595 12733
rect 4065 12699 4123 12705
rect 4065 12665 4077 12699
rect 4111 12665 4123 12699
rect 4065 12659 4123 12665
rect 4709 12699 4767 12705
rect 4709 12665 4721 12699
rect 4755 12696 4767 12699
rect 4798 12696 4804 12708
rect 4755 12668 4804 12696
rect 4755 12665 4767 12668
rect 4709 12659 4767 12665
rect 1670 12628 1676 12640
rect 1631 12600 1676 12628
rect 1670 12588 1676 12600
rect 1728 12588 1734 12640
rect 2130 12628 2136 12640
rect 2091 12600 2136 12628
rect 2130 12588 2136 12600
rect 2188 12588 2194 12640
rect 4080 12628 4108 12659
rect 4798 12656 4804 12668
rect 4856 12656 4862 12708
rect 4893 12699 4951 12705
rect 4893 12665 4905 12699
rect 4939 12696 4951 12699
rect 5350 12696 5356 12708
rect 4939 12668 5356 12696
rect 4939 12665 4951 12668
rect 4893 12659 4951 12665
rect 5350 12656 5356 12668
rect 5408 12656 5414 12708
rect 5445 12699 5503 12705
rect 5445 12665 5457 12699
rect 5491 12696 5503 12699
rect 6270 12696 6276 12708
rect 5491 12668 6276 12696
rect 5491 12665 5503 12668
rect 5445 12659 5503 12665
rect 6270 12656 6276 12668
rect 6328 12656 6334 12708
rect 6914 12696 6920 12708
rect 6875 12668 6920 12696
rect 6914 12656 6920 12668
rect 6972 12656 6978 12708
rect 7392 12696 7420 12804
rect 8846 12792 8852 12804
rect 8904 12792 8910 12844
rect 7466 12724 7472 12776
rect 7524 12764 7530 12776
rect 7653 12767 7711 12773
rect 7653 12764 7665 12767
rect 7524 12736 7665 12764
rect 7524 12724 7530 12736
rect 7653 12733 7665 12736
rect 7699 12733 7711 12767
rect 7653 12727 7711 12733
rect 7742 12724 7748 12776
rect 7800 12764 7806 12776
rect 8297 12767 8355 12773
rect 8297 12764 8309 12767
rect 7800 12736 8309 12764
rect 7800 12724 7806 12736
rect 8297 12733 8309 12736
rect 8343 12764 8355 12767
rect 8956 12764 8984 12872
rect 9493 12869 9505 12903
rect 9539 12900 9551 12903
rect 10870 12900 10876 12912
rect 9539 12872 10876 12900
rect 9539 12869 9551 12872
rect 9493 12863 9551 12869
rect 10870 12860 10876 12872
rect 10928 12860 10934 12912
rect 9033 12835 9091 12841
rect 9033 12801 9045 12835
rect 9079 12832 9091 12835
rect 9858 12832 9864 12844
rect 9079 12804 9864 12832
rect 9079 12801 9091 12804
rect 9033 12795 9091 12801
rect 9858 12792 9864 12804
rect 9916 12792 9922 12844
rect 10226 12832 10232 12844
rect 10187 12804 10232 12832
rect 10226 12792 10232 12804
rect 10284 12792 10290 12844
rect 10410 12832 10416 12844
rect 10371 12804 10416 12832
rect 10410 12792 10416 12804
rect 10468 12792 10474 12844
rect 11238 12792 11244 12844
rect 11296 12832 11302 12844
rect 11333 12835 11391 12841
rect 11333 12832 11345 12835
rect 11296 12804 11345 12832
rect 11296 12792 11302 12804
rect 11333 12801 11345 12804
rect 11379 12801 11391 12835
rect 11333 12795 11391 12801
rect 10137 12767 10195 12773
rect 10137 12764 10149 12767
rect 8343 12736 8892 12764
rect 8956 12736 10149 12764
rect 8343 12733 8355 12736
rect 8297 12727 8355 12733
rect 8864 12708 8892 12736
rect 10137 12733 10149 12736
rect 10183 12733 10195 12767
rect 10137 12727 10195 12733
rect 10781 12767 10839 12773
rect 10781 12733 10793 12767
rect 10827 12764 10839 12767
rect 11701 12767 11759 12773
rect 11701 12764 11713 12767
rect 10827 12736 11713 12764
rect 10827 12733 10839 12736
rect 10781 12727 10839 12733
rect 11701 12733 11713 12736
rect 11747 12764 11759 12767
rect 11790 12764 11796 12776
rect 11747 12736 11796 12764
rect 11747 12733 11759 12736
rect 11701 12727 11759 12733
rect 11790 12724 11796 12736
rect 11848 12724 11854 12776
rect 13170 12764 13176 12776
rect 13131 12736 13176 12764
rect 13170 12724 13176 12736
rect 13228 12724 13234 12776
rect 7926 12696 7932 12708
rect 7392 12668 7932 12696
rect 7926 12656 7932 12668
rect 7984 12656 7990 12708
rect 8018 12656 8024 12708
rect 8076 12696 8082 12708
rect 8481 12699 8539 12705
rect 8481 12696 8493 12699
rect 8076 12668 8493 12696
rect 8076 12656 8082 12668
rect 8481 12665 8493 12668
rect 8527 12696 8539 12699
rect 8662 12696 8668 12708
rect 8527 12668 8668 12696
rect 8527 12665 8539 12668
rect 8481 12659 8539 12665
rect 8662 12656 8668 12668
rect 8720 12656 8726 12708
rect 8846 12656 8852 12708
rect 8904 12656 8910 12708
rect 11241 12699 11299 12705
rect 11241 12665 11253 12699
rect 11287 12696 11299 12699
rect 11882 12696 11888 12708
rect 11287 12668 11888 12696
rect 11287 12665 11299 12668
rect 11241 12659 11299 12665
rect 11882 12656 11888 12668
rect 11940 12696 11946 12708
rect 13265 12699 13323 12705
rect 13265 12696 13277 12699
rect 11940 12668 13277 12696
rect 11940 12656 11946 12668
rect 13265 12665 13277 12668
rect 13311 12665 13323 12699
rect 13265 12659 13323 12665
rect 5994 12628 6000 12640
rect 4080 12600 6000 12628
rect 5994 12588 6000 12600
rect 6052 12588 6058 12640
rect 7006 12628 7012 12640
rect 6967 12600 7012 12628
rect 7006 12588 7012 12600
rect 7064 12588 7070 12640
rect 7374 12628 7380 12640
rect 7335 12600 7380 12628
rect 7374 12588 7380 12600
rect 7432 12588 7438 12640
rect 7745 12631 7803 12637
rect 7745 12597 7757 12631
rect 7791 12628 7803 12631
rect 8570 12628 8576 12640
rect 7791 12600 8576 12628
rect 7791 12597 7803 12600
rect 7745 12591 7803 12597
rect 8570 12588 8576 12600
rect 8628 12588 8634 12640
rect 9125 12631 9183 12637
rect 9125 12597 9137 12631
rect 9171 12628 9183 12631
rect 9214 12628 9220 12640
rect 9171 12600 9220 12628
rect 9171 12597 9183 12600
rect 9125 12591 9183 12597
rect 9214 12588 9220 12600
rect 9272 12588 9278 12640
rect 1104 12538 13892 12560
rect 1104 12486 8246 12538
rect 8298 12486 8310 12538
rect 8362 12486 8374 12538
rect 8426 12486 8438 12538
rect 8490 12486 13892 12538
rect 1104 12464 13892 12486
rect 4338 12424 4344 12436
rect 4299 12396 4344 12424
rect 4338 12384 4344 12396
rect 4396 12384 4402 12436
rect 5534 12384 5540 12436
rect 5592 12424 5598 12436
rect 5905 12427 5963 12433
rect 5905 12424 5917 12427
rect 5592 12396 5917 12424
rect 5592 12384 5598 12396
rect 5905 12393 5917 12396
rect 5951 12393 5963 12427
rect 5905 12387 5963 12393
rect 7006 12384 7012 12436
rect 7064 12424 7070 12436
rect 7190 12424 7196 12436
rect 7064 12396 7196 12424
rect 7064 12384 7070 12396
rect 7190 12384 7196 12396
rect 7248 12424 7254 12436
rect 7285 12427 7343 12433
rect 7285 12424 7297 12427
rect 7248 12396 7297 12424
rect 7248 12384 7254 12396
rect 7285 12393 7297 12396
rect 7331 12393 7343 12427
rect 9122 12424 9128 12436
rect 7285 12387 7343 12393
rect 7392 12396 9128 12424
rect 3050 12356 3056 12368
rect 3011 12328 3056 12356
rect 3050 12316 3056 12328
rect 3108 12316 3114 12368
rect 4798 12316 4804 12368
rect 4856 12356 4862 12368
rect 5258 12356 5264 12368
rect 4856 12328 5264 12356
rect 4856 12316 4862 12328
rect 5258 12316 5264 12328
rect 5316 12316 5322 12368
rect 7392 12356 7420 12396
rect 9122 12384 9128 12396
rect 9180 12384 9186 12436
rect 9306 12424 9312 12436
rect 9267 12396 9312 12424
rect 9306 12384 9312 12396
rect 9364 12384 9370 12436
rect 9769 12427 9827 12433
rect 9769 12393 9781 12427
rect 9815 12424 9827 12427
rect 10318 12424 10324 12436
rect 9815 12396 10324 12424
rect 9815 12393 9827 12396
rect 9769 12387 9827 12393
rect 10318 12384 10324 12396
rect 10376 12384 10382 12436
rect 11422 12384 11428 12436
rect 11480 12424 11486 12436
rect 12345 12427 12403 12433
rect 12345 12424 12357 12427
rect 11480 12396 12357 12424
rect 11480 12384 11486 12396
rect 12345 12393 12357 12396
rect 12391 12393 12403 12427
rect 12345 12387 12403 12393
rect 13081 12427 13139 12433
rect 13081 12393 13093 12427
rect 13127 12424 13139 12427
rect 13170 12424 13176 12436
rect 13127 12396 13176 12424
rect 13127 12393 13139 12396
rect 13081 12387 13139 12393
rect 13170 12384 13176 12396
rect 13228 12384 13234 12436
rect 5460 12328 7420 12356
rect 1489 12291 1547 12297
rect 1489 12257 1501 12291
rect 1535 12288 1547 12291
rect 2130 12288 2136 12300
rect 1535 12260 2136 12288
rect 1535 12257 1547 12260
rect 1489 12251 1547 12257
rect 2130 12248 2136 12260
rect 2188 12248 2194 12300
rect 2774 12248 2780 12300
rect 2832 12288 2838 12300
rect 3329 12291 3387 12297
rect 2832 12260 2877 12288
rect 2832 12248 2838 12260
rect 3329 12257 3341 12291
rect 3375 12288 3387 12291
rect 4062 12288 4068 12300
rect 3375 12260 4068 12288
rect 3375 12257 3387 12260
rect 3329 12251 3387 12257
rect 4062 12248 4068 12260
rect 4120 12248 4126 12300
rect 4249 12291 4307 12297
rect 4249 12257 4261 12291
rect 4295 12288 4307 12291
rect 4893 12291 4951 12297
rect 4893 12288 4905 12291
rect 4295 12260 4905 12288
rect 4295 12257 4307 12260
rect 4249 12251 4307 12257
rect 4893 12257 4905 12260
rect 4939 12257 4951 12291
rect 5166 12288 5172 12300
rect 5127 12260 5172 12288
rect 4893 12251 4951 12257
rect 5166 12248 5172 12260
rect 5224 12248 5230 12300
rect 2038 12180 2044 12232
rect 2096 12220 2102 12232
rect 4525 12223 4583 12229
rect 4525 12220 4537 12223
rect 2096 12192 4537 12220
rect 2096 12180 2102 12192
rect 4525 12189 4537 12192
rect 4571 12189 4583 12223
rect 5276 12220 5304 12316
rect 5460 12300 5488 12328
rect 5442 12288 5448 12300
rect 5355 12260 5448 12288
rect 5442 12248 5448 12260
rect 5500 12248 5506 12300
rect 6380 12297 6408 12328
rect 7558 12316 7564 12368
rect 7616 12356 7622 12368
rect 7616 12328 8524 12356
rect 7616 12316 7622 12328
rect 8496 12300 8524 12328
rect 9490 12316 9496 12368
rect 9548 12356 9554 12368
rect 10226 12356 10232 12368
rect 9548 12328 10232 12356
rect 9548 12316 9554 12328
rect 10226 12316 10232 12328
rect 10284 12356 10290 12368
rect 11698 12356 11704 12368
rect 10284 12328 10364 12356
rect 11659 12328 11704 12356
rect 10284 12316 10290 12328
rect 5721 12291 5779 12297
rect 5721 12257 5733 12291
rect 5767 12288 5779 12291
rect 6089 12291 6147 12297
rect 6089 12288 6101 12291
rect 5767 12260 6101 12288
rect 5767 12257 5779 12260
rect 5721 12251 5779 12257
rect 6089 12257 6101 12260
rect 6135 12257 6147 12291
rect 6089 12251 6147 12257
rect 6365 12291 6423 12297
rect 6365 12257 6377 12291
rect 6411 12257 6423 12291
rect 6365 12251 6423 12257
rect 6733 12291 6791 12297
rect 6733 12257 6745 12291
rect 6779 12288 6791 12291
rect 7374 12288 7380 12300
rect 6779 12260 7380 12288
rect 6779 12257 6791 12260
rect 6733 12251 6791 12257
rect 5353 12223 5411 12229
rect 5353 12220 5365 12223
rect 5276 12192 5365 12220
rect 4525 12183 4583 12189
rect 5353 12189 5365 12192
rect 5399 12220 5411 12223
rect 6748 12220 6776 12251
rect 7374 12248 7380 12260
rect 7432 12288 7438 12300
rect 7469 12291 7527 12297
rect 7469 12288 7481 12291
rect 7432 12260 7481 12288
rect 7432 12248 7438 12260
rect 7469 12257 7481 12260
rect 7515 12257 7527 12291
rect 7742 12288 7748 12300
rect 7703 12260 7748 12288
rect 7469 12251 7527 12257
rect 7742 12248 7748 12260
rect 7800 12248 7806 12300
rect 7929 12291 7987 12297
rect 7929 12257 7941 12291
rect 7975 12288 7987 12291
rect 8018 12288 8024 12300
rect 7975 12260 8024 12288
rect 7975 12257 7987 12260
rect 7929 12251 7987 12257
rect 8018 12248 8024 12260
rect 8076 12248 8082 12300
rect 8478 12288 8484 12300
rect 8391 12260 8484 12288
rect 8478 12248 8484 12260
rect 8536 12248 8542 12300
rect 8665 12291 8723 12297
rect 8665 12257 8677 12291
rect 8711 12288 8723 12291
rect 8754 12288 8760 12300
rect 8711 12260 8760 12288
rect 8711 12257 8723 12260
rect 8665 12251 8723 12257
rect 8754 12248 8760 12260
rect 8812 12248 8818 12300
rect 9677 12291 9735 12297
rect 9677 12257 9689 12291
rect 9723 12288 9735 12291
rect 10134 12288 10140 12300
rect 9723 12260 10140 12288
rect 9723 12257 9735 12260
rect 9677 12251 9735 12257
rect 10134 12248 10140 12260
rect 10192 12248 10198 12300
rect 10336 12297 10364 12328
rect 11698 12316 11704 12328
rect 11756 12316 11762 12368
rect 10321 12291 10379 12297
rect 10321 12257 10333 12291
rect 10367 12257 10379 12291
rect 10321 12251 10379 12257
rect 10505 12291 10563 12297
rect 10505 12257 10517 12291
rect 10551 12288 10563 12291
rect 10594 12288 10600 12300
rect 10551 12260 10600 12288
rect 10551 12257 10563 12260
rect 10505 12251 10563 12257
rect 10594 12248 10600 12260
rect 10652 12248 10658 12300
rect 11149 12291 11207 12297
rect 11149 12257 11161 12291
rect 11195 12288 11207 12291
rect 11330 12288 11336 12300
rect 11195 12260 11336 12288
rect 11195 12257 11207 12260
rect 11149 12251 11207 12257
rect 11330 12248 11336 12260
rect 11388 12248 11394 12300
rect 11606 12288 11612 12300
rect 11567 12260 11612 12288
rect 11606 12248 11612 12260
rect 11664 12248 11670 12300
rect 13170 12288 13176 12300
rect 13131 12260 13176 12288
rect 13170 12248 13176 12260
rect 13228 12248 13234 12300
rect 5399 12192 6776 12220
rect 5399 12189 5411 12192
rect 5353 12183 5411 12189
rect 3142 12112 3148 12164
rect 3200 12152 3206 12164
rect 3881 12155 3939 12161
rect 3881 12152 3893 12155
rect 3200 12124 3893 12152
rect 3200 12112 3206 12124
rect 3881 12121 3893 12124
rect 3927 12121 3939 12155
rect 4540 12152 4568 12183
rect 6822 12180 6828 12232
rect 6880 12220 6886 12232
rect 7653 12223 7711 12229
rect 7653 12220 7665 12223
rect 6880 12192 7665 12220
rect 6880 12180 6886 12192
rect 7653 12189 7665 12192
rect 7699 12220 7711 12223
rect 8110 12220 8116 12232
rect 7699 12192 8116 12220
rect 7699 12189 7711 12192
rect 7653 12183 7711 12189
rect 8110 12180 8116 12192
rect 8168 12220 8174 12232
rect 8386 12220 8392 12232
rect 8168 12192 8392 12220
rect 8168 12180 8174 12192
rect 8386 12180 8392 12192
rect 8444 12180 8450 12232
rect 9953 12223 10011 12229
rect 9953 12189 9965 12223
rect 9999 12189 10011 12223
rect 9953 12183 10011 12189
rect 4890 12152 4896 12164
rect 4540 12124 4896 12152
rect 3881 12115 3939 12121
rect 4890 12112 4896 12124
rect 4948 12112 4954 12164
rect 5265 12155 5323 12161
rect 5265 12121 5277 12155
rect 5311 12152 5323 12155
rect 6086 12152 6092 12164
rect 5311 12124 6092 12152
rect 5311 12121 5323 12124
rect 5265 12115 5323 12121
rect 6086 12112 6092 12124
rect 6144 12152 6150 12164
rect 6185 12155 6243 12161
rect 6185 12152 6197 12155
rect 6144 12124 6197 12152
rect 6144 12112 6150 12124
rect 6185 12121 6197 12124
rect 6231 12121 6243 12155
rect 6185 12115 6243 12121
rect 6273 12155 6331 12161
rect 6273 12121 6285 12155
rect 6319 12121 6331 12155
rect 6273 12115 6331 12121
rect 3513 12087 3571 12093
rect 3513 12053 3525 12087
rect 3559 12084 3571 12087
rect 3786 12084 3792 12096
rect 3559 12056 3792 12084
rect 3559 12053 3571 12056
rect 3513 12047 3571 12053
rect 3786 12044 3792 12056
rect 3844 12044 3850 12096
rect 5166 12044 5172 12096
rect 5224 12084 5230 12096
rect 5626 12084 5632 12096
rect 5224 12056 5632 12084
rect 5224 12044 5230 12056
rect 5626 12044 5632 12056
rect 5684 12084 5690 12096
rect 5721 12087 5779 12093
rect 5721 12084 5733 12087
rect 5684 12056 5733 12084
rect 5684 12044 5690 12056
rect 5721 12053 5733 12056
rect 5767 12053 5779 12087
rect 6288 12084 6316 12115
rect 7282 12112 7288 12164
rect 7340 12152 7346 12164
rect 7561 12155 7619 12161
rect 7561 12152 7573 12155
rect 7340 12124 7573 12152
rect 7340 12112 7346 12124
rect 7561 12121 7573 12124
rect 7607 12121 7619 12155
rect 9968 12152 9996 12183
rect 12066 12180 12072 12232
rect 12124 12220 12130 12232
rect 12437 12223 12495 12229
rect 12437 12220 12449 12223
rect 12124 12192 12449 12220
rect 12124 12180 12130 12192
rect 12437 12189 12449 12192
rect 12483 12189 12495 12223
rect 12437 12183 12495 12189
rect 12529 12223 12587 12229
rect 12529 12189 12541 12223
rect 12575 12220 12587 12223
rect 12575 12192 12609 12220
rect 12575 12189 12587 12192
rect 12529 12183 12587 12189
rect 10410 12152 10416 12164
rect 9968 12124 10416 12152
rect 7561 12115 7619 12121
rect 10410 12112 10416 12124
rect 10468 12152 10474 12164
rect 12544 12152 12572 12183
rect 12802 12152 12808 12164
rect 10468 12124 12808 12152
rect 10468 12112 10474 12124
rect 12802 12112 12808 12124
rect 12860 12112 12866 12164
rect 6362 12084 6368 12096
rect 6288 12056 6368 12084
rect 5721 12047 5779 12053
rect 6362 12044 6368 12056
rect 6420 12044 6426 12096
rect 6825 12087 6883 12093
rect 6825 12053 6837 12087
rect 6871 12084 6883 12087
rect 6914 12084 6920 12096
rect 6871 12056 6920 12084
rect 6871 12053 6883 12056
rect 6825 12047 6883 12053
rect 6914 12044 6920 12056
rect 6972 12044 6978 12096
rect 7006 12044 7012 12096
rect 7064 12084 7070 12096
rect 8297 12087 8355 12093
rect 8297 12084 8309 12087
rect 7064 12056 8309 12084
rect 7064 12044 7070 12056
rect 8297 12053 8309 12056
rect 8343 12053 8355 12087
rect 8478 12084 8484 12096
rect 8439 12056 8484 12084
rect 8297 12047 8355 12053
rect 8478 12044 8484 12056
rect 8536 12044 8542 12096
rect 9306 12044 9312 12096
rect 9364 12084 9370 12096
rect 10597 12087 10655 12093
rect 10597 12084 10609 12087
rect 9364 12056 10609 12084
rect 9364 12044 9370 12056
rect 10597 12053 10609 12056
rect 10643 12053 10655 12087
rect 11974 12084 11980 12096
rect 11935 12056 11980 12084
rect 10597 12047 10655 12053
rect 11974 12044 11980 12056
rect 12032 12044 12038 12096
rect 1104 11994 13892 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 12246 11994
rect 12298 11942 12310 11994
rect 12362 11942 12374 11994
rect 12426 11942 12438 11994
rect 12490 11942 13892 11994
rect 1104 11920 13892 11942
rect 5994 11880 6000 11892
rect 5955 11852 6000 11880
rect 5994 11840 6000 11852
rect 6052 11840 6058 11892
rect 6546 11880 6552 11892
rect 6507 11852 6552 11880
rect 6546 11840 6552 11852
rect 6604 11840 6610 11892
rect 8478 11880 8484 11892
rect 7024 11852 8484 11880
rect 5074 11812 5080 11824
rect 5035 11784 5080 11812
rect 5074 11772 5080 11784
rect 5132 11772 5138 11824
rect 6730 11772 6736 11824
rect 6788 11812 6794 11824
rect 6917 11815 6975 11821
rect 6917 11812 6929 11815
rect 6788 11784 6929 11812
rect 6788 11772 6794 11784
rect 6917 11781 6929 11784
rect 6963 11781 6975 11815
rect 6917 11775 6975 11781
rect 474 11704 480 11756
rect 532 11744 538 11756
rect 2225 11747 2283 11753
rect 2225 11744 2237 11747
rect 532 11716 2237 11744
rect 532 11704 538 11716
rect 2225 11713 2237 11716
rect 2271 11713 2283 11747
rect 2225 11707 2283 11713
rect 2317 11747 2375 11753
rect 2317 11713 2329 11747
rect 2363 11713 2375 11747
rect 5534 11744 5540 11756
rect 2317 11707 2375 11713
rect 3896 11716 5540 11744
rect 2038 11636 2044 11688
rect 2096 11676 2102 11688
rect 2332 11676 2360 11707
rect 3142 11676 3148 11688
rect 2096 11648 2360 11676
rect 3103 11648 3148 11676
rect 2096 11636 2102 11648
rect 3142 11636 3148 11648
rect 3200 11636 3206 11688
rect 3418 11676 3424 11688
rect 3379 11648 3424 11676
rect 3418 11636 3424 11648
rect 3476 11636 3482 11688
rect 2133 11611 2191 11617
rect 2133 11577 2145 11611
rect 2179 11608 2191 11611
rect 2179 11580 2452 11608
rect 2179 11577 2191 11580
rect 2133 11571 2191 11577
rect 1762 11540 1768 11552
rect 1723 11512 1768 11540
rect 1762 11500 1768 11512
rect 1820 11500 1826 11552
rect 2424 11540 2452 11580
rect 2774 11568 2780 11620
rect 2832 11608 2838 11620
rect 2961 11611 3019 11617
rect 2832 11580 2877 11608
rect 2832 11568 2838 11580
rect 2961 11577 2973 11611
rect 3007 11608 3019 11611
rect 3326 11608 3332 11620
rect 3007 11580 3332 11608
rect 3007 11577 3019 11580
rect 2961 11571 3019 11577
rect 3326 11568 3332 11580
rect 3384 11568 3390 11620
rect 3896 11540 3924 11716
rect 5534 11704 5540 11716
rect 5592 11704 5598 11756
rect 6086 11704 6092 11756
rect 6144 11744 6150 11756
rect 7024 11753 7052 11852
rect 8478 11840 8484 11852
rect 8536 11840 8542 11892
rect 10134 11840 10140 11892
rect 10192 11880 10198 11892
rect 11701 11883 11759 11889
rect 10192 11852 10916 11880
rect 10192 11840 10198 11852
rect 8297 11815 8355 11821
rect 8297 11781 8309 11815
rect 8343 11812 8355 11815
rect 8570 11812 8576 11824
rect 8343 11784 8576 11812
rect 8343 11781 8355 11784
rect 8297 11775 8355 11781
rect 8570 11772 8576 11784
rect 8628 11772 8634 11824
rect 9214 11772 9220 11824
rect 9272 11812 9278 11824
rect 10888 11821 10916 11852
rect 11701 11849 11713 11883
rect 11747 11880 11759 11883
rect 11790 11880 11796 11892
rect 11747 11852 11796 11880
rect 11747 11849 11759 11852
rect 11701 11843 11759 11849
rect 11790 11840 11796 11852
rect 11848 11840 11854 11892
rect 9489 11815 9547 11821
rect 9489 11812 9501 11815
rect 9272 11784 9501 11812
rect 9272 11772 9278 11784
rect 9489 11781 9501 11784
rect 9535 11781 9547 11815
rect 9489 11775 9547 11781
rect 10873 11815 10931 11821
rect 10873 11781 10885 11815
rect 10919 11781 10931 11815
rect 13170 11812 13176 11824
rect 13131 11784 13176 11812
rect 10873 11775 10931 11781
rect 13170 11772 13176 11784
rect 13228 11772 13234 11824
rect 7009 11747 7067 11753
rect 7009 11744 7021 11747
rect 6144 11716 7021 11744
rect 6144 11704 6150 11716
rect 7009 11713 7021 11716
rect 7055 11713 7067 11747
rect 7009 11707 7067 11713
rect 7101 11747 7159 11753
rect 7101 11713 7113 11747
rect 7147 11744 7159 11747
rect 7282 11744 7288 11756
rect 7147 11716 7288 11744
rect 7147 11713 7159 11716
rect 7101 11707 7159 11713
rect 7282 11704 7288 11716
rect 7340 11704 7346 11756
rect 8386 11744 8392 11756
rect 8347 11716 8392 11744
rect 8386 11704 8392 11716
rect 8444 11704 8450 11756
rect 8846 11744 8852 11756
rect 8496 11716 8852 11744
rect 3970 11636 3976 11688
rect 4028 11676 4034 11688
rect 4157 11679 4215 11685
rect 4157 11676 4169 11679
rect 4028 11648 4169 11676
rect 4028 11636 4034 11648
rect 4157 11645 4169 11648
rect 4203 11676 4215 11679
rect 5905 11679 5963 11685
rect 5905 11676 5917 11679
rect 4203 11648 5917 11676
rect 4203 11645 4215 11648
rect 4157 11639 4215 11645
rect 5905 11645 5917 11648
rect 5951 11645 5963 11679
rect 5905 11639 5963 11645
rect 6454 11636 6460 11688
rect 6512 11676 6518 11688
rect 6825 11679 6883 11685
rect 6825 11676 6837 11679
rect 6512 11648 6837 11676
rect 6512 11636 6518 11648
rect 6825 11645 6837 11648
rect 6871 11645 6883 11679
rect 6825 11639 6883 11645
rect 7193 11679 7251 11685
rect 7193 11645 7205 11679
rect 7239 11676 7251 11679
rect 7374 11676 7380 11688
rect 7239 11648 7380 11676
rect 7239 11645 7251 11648
rect 7193 11639 7251 11645
rect 7374 11636 7380 11648
rect 7432 11636 7438 11688
rect 8018 11676 8024 11688
rect 7979 11648 8024 11676
rect 8018 11636 8024 11648
rect 8076 11636 8082 11688
rect 8496 11685 8524 11716
rect 8846 11704 8852 11716
rect 8904 11744 8910 11756
rect 9122 11744 9128 11756
rect 8904 11716 9128 11744
rect 8904 11704 8910 11716
rect 9122 11704 9128 11716
rect 9180 11744 9186 11756
rect 9401 11747 9459 11753
rect 9401 11744 9413 11747
rect 9180 11716 9413 11744
rect 9180 11704 9186 11716
rect 9401 11713 9413 11716
rect 9447 11713 9459 11747
rect 9401 11707 9459 11713
rect 9674 11704 9680 11756
rect 9732 11744 9738 11756
rect 10502 11744 10508 11756
rect 9732 11716 10508 11744
rect 9732 11704 9738 11716
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 12345 11747 12403 11753
rect 12345 11713 12357 11747
rect 12391 11744 12403 11747
rect 12802 11744 12808 11756
rect 12391 11716 12808 11744
rect 12391 11713 12403 11716
rect 12345 11707 12403 11713
rect 12802 11704 12808 11716
rect 12860 11704 12866 11756
rect 13262 11744 13268 11756
rect 13223 11716 13268 11744
rect 13262 11704 13268 11716
rect 13320 11704 13326 11756
rect 8205 11679 8263 11685
rect 8205 11676 8217 11679
rect 8128 11648 8217 11676
rect 8128 11620 8156 11648
rect 8205 11645 8217 11648
rect 8251 11645 8263 11679
rect 8205 11639 8263 11645
rect 8481 11679 8539 11685
rect 8481 11645 8493 11679
rect 8527 11645 8539 11679
rect 8662 11676 8668 11688
rect 8575 11648 8668 11676
rect 8481 11639 8539 11645
rect 8662 11636 8668 11648
rect 8720 11636 8726 11688
rect 9306 11676 9312 11688
rect 9267 11648 9312 11676
rect 9306 11636 9312 11648
rect 9364 11636 9370 11688
rect 9585 11679 9643 11685
rect 9585 11645 9597 11679
rect 9631 11645 9643 11679
rect 9585 11639 9643 11645
rect 9861 11679 9919 11685
rect 9861 11645 9873 11679
rect 9907 11676 9919 11679
rect 10962 11676 10968 11688
rect 9907 11648 10824 11676
rect 10923 11648 10968 11676
rect 9907 11645 9919 11648
rect 9861 11639 9919 11645
rect 4062 11568 4068 11620
rect 4120 11608 4126 11620
rect 4341 11611 4399 11617
rect 4341 11608 4353 11611
rect 4120 11580 4353 11608
rect 4120 11568 4126 11580
rect 4341 11577 4353 11580
rect 4387 11577 4399 11611
rect 5258 11608 5264 11620
rect 5219 11580 5264 11608
rect 4341 11571 4399 11577
rect 5258 11568 5264 11580
rect 5316 11568 5322 11620
rect 5626 11608 5632 11620
rect 5587 11580 5632 11608
rect 5626 11568 5632 11580
rect 5684 11568 5690 11620
rect 6362 11568 6368 11620
rect 6420 11608 6426 11620
rect 8110 11608 8116 11620
rect 6420 11580 8116 11608
rect 6420 11568 6426 11580
rect 8110 11568 8116 11580
rect 8168 11568 8174 11620
rect 8680 11608 8708 11636
rect 9398 11608 9404 11620
rect 8680 11580 9404 11608
rect 9398 11568 9404 11580
rect 9456 11568 9462 11620
rect 9600 11608 9628 11639
rect 10137 11611 10195 11617
rect 9600 11580 9904 11608
rect 9876 11552 9904 11580
rect 10137 11577 10149 11611
rect 10183 11608 10195 11611
rect 10226 11608 10232 11620
rect 10183 11580 10232 11608
rect 10183 11577 10195 11580
rect 10137 11571 10195 11577
rect 10226 11568 10232 11580
rect 10284 11568 10290 11620
rect 10321 11611 10379 11617
rect 10321 11577 10333 11611
rect 10367 11577 10379 11611
rect 10796 11608 10824 11648
rect 10962 11636 10968 11648
rect 11020 11636 11026 11688
rect 11149 11679 11207 11685
rect 11149 11645 11161 11679
rect 11195 11676 11207 11679
rect 11790 11676 11796 11688
rect 11195 11648 11796 11676
rect 11195 11645 11207 11648
rect 11149 11639 11207 11645
rect 11790 11636 11796 11648
rect 11848 11636 11854 11688
rect 11974 11636 11980 11688
rect 12032 11676 12038 11688
rect 12713 11679 12771 11685
rect 12713 11676 12725 11679
rect 12032 11648 12725 11676
rect 12032 11636 12038 11648
rect 12713 11645 12725 11648
rect 12759 11645 12771 11679
rect 12713 11639 12771 11645
rect 12069 11611 12127 11617
rect 12069 11608 12081 11611
rect 10796 11580 12081 11608
rect 10321 11571 10379 11577
rect 12069 11577 12081 11580
rect 12115 11577 12127 11611
rect 12069 11571 12127 11577
rect 2424 11512 3924 11540
rect 4617 11543 4675 11549
rect 4617 11509 4629 11543
rect 4663 11540 4675 11543
rect 4706 11540 4712 11552
rect 4663 11512 4712 11540
rect 4663 11509 4675 11512
rect 4617 11503 4675 11509
rect 4706 11500 4712 11512
rect 4764 11500 4770 11552
rect 5350 11540 5356 11552
rect 5311 11512 5356 11540
rect 5350 11500 5356 11512
rect 5408 11500 5414 11552
rect 5445 11543 5503 11549
rect 5445 11509 5457 11543
rect 5491 11540 5503 11543
rect 5718 11540 5724 11552
rect 5491 11512 5724 11540
rect 5491 11509 5503 11512
rect 5445 11503 5503 11509
rect 5718 11500 5724 11512
rect 5776 11500 5782 11552
rect 5902 11500 5908 11552
rect 5960 11540 5966 11552
rect 8662 11540 8668 11552
rect 5960 11512 8668 11540
rect 5960 11500 5966 11512
rect 8662 11500 8668 11512
rect 8720 11500 8726 11552
rect 9858 11500 9864 11552
rect 9916 11540 9922 11552
rect 10336 11540 10364 11571
rect 9916 11512 10364 11540
rect 9916 11500 9922 11512
rect 11882 11500 11888 11552
rect 11940 11540 11946 11552
rect 12161 11543 12219 11549
rect 12161 11540 12173 11543
rect 11940 11512 12173 11540
rect 11940 11500 11946 11512
rect 12161 11509 12173 11512
rect 12207 11509 12219 11543
rect 12161 11503 12219 11509
rect 1104 11450 13892 11472
rect 1104 11398 8246 11450
rect 8298 11398 8310 11450
rect 8362 11398 8374 11450
rect 8426 11398 8438 11450
rect 8490 11398 13892 11450
rect 1104 11376 13892 11398
rect 3418 11296 3424 11348
rect 3476 11336 3482 11348
rect 7653 11339 7711 11345
rect 7653 11336 7665 11339
rect 3476 11308 7665 11336
rect 3476 11296 3482 11308
rect 1780 11240 3556 11268
rect 1780 11212 1808 11240
rect 1762 11200 1768 11212
rect 1723 11172 1768 11200
rect 1762 11160 1768 11172
rect 1820 11160 1826 11212
rect 2406 11200 2412 11212
rect 2367 11172 2412 11200
rect 2406 11160 2412 11172
rect 2464 11160 2470 11212
rect 2682 11200 2688 11212
rect 2643 11172 2688 11200
rect 2682 11160 2688 11172
rect 2740 11160 2746 11212
rect 3528 11209 3556 11240
rect 3786 11228 3792 11280
rect 3844 11268 3850 11280
rect 3881 11271 3939 11277
rect 3881 11268 3893 11271
rect 3844 11240 3893 11268
rect 3844 11228 3850 11240
rect 3881 11237 3893 11240
rect 3927 11237 3939 11271
rect 3881 11231 3939 11237
rect 3970 11228 3976 11280
rect 4028 11268 4034 11280
rect 4028 11240 4073 11268
rect 4028 11228 4034 11240
rect 4448 11209 4476 11308
rect 7653 11305 7665 11308
rect 7699 11305 7711 11339
rect 8018 11336 8024 11348
rect 7979 11308 8024 11336
rect 7653 11299 7711 11305
rect 8018 11296 8024 11308
rect 8076 11296 8082 11348
rect 9585 11339 9643 11345
rect 9585 11305 9597 11339
rect 9631 11336 9643 11339
rect 9766 11336 9772 11348
rect 9631 11308 9772 11336
rect 9631 11305 9643 11308
rect 9585 11299 9643 11305
rect 9766 11296 9772 11308
rect 9824 11296 9830 11348
rect 10502 11296 10508 11348
rect 10560 11336 10566 11348
rect 11057 11339 11115 11345
rect 11057 11336 11069 11339
rect 10560 11308 11069 11336
rect 10560 11296 10566 11308
rect 11057 11305 11069 11308
rect 11103 11305 11115 11339
rect 11057 11299 11115 11305
rect 5629 11271 5687 11277
rect 5629 11237 5641 11271
rect 5675 11268 5687 11271
rect 5902 11268 5908 11280
rect 5675 11240 5908 11268
rect 5675 11237 5687 11240
rect 5629 11231 5687 11237
rect 5902 11228 5908 11240
rect 5960 11228 5966 11280
rect 6089 11271 6147 11277
rect 6089 11237 6101 11271
rect 6135 11268 6147 11271
rect 7834 11268 7840 11280
rect 6135 11240 7840 11268
rect 6135 11237 6147 11240
rect 6089 11231 6147 11237
rect 7834 11228 7840 11240
rect 7892 11228 7898 11280
rect 8113 11271 8171 11277
rect 8113 11237 8125 11271
rect 8159 11268 8171 11271
rect 9030 11268 9036 11280
rect 8159 11240 9036 11268
rect 8159 11237 8171 11240
rect 8113 11231 8171 11237
rect 9030 11228 9036 11240
rect 9088 11228 9094 11280
rect 10042 11228 10048 11280
rect 10100 11268 10106 11280
rect 10962 11268 10968 11280
rect 10100 11240 10968 11268
rect 10100 11228 10106 11240
rect 10962 11228 10968 11240
rect 11020 11228 11026 11280
rect 13170 11228 13176 11280
rect 13228 11268 13234 11280
rect 13357 11271 13415 11277
rect 13357 11268 13369 11271
rect 13228 11240 13369 11268
rect 13228 11228 13234 11240
rect 13357 11237 13369 11240
rect 13403 11237 13415 11271
rect 13357 11231 13415 11237
rect 3513 11203 3571 11209
rect 3513 11169 3525 11203
rect 3559 11169 3571 11203
rect 3513 11163 3571 11169
rect 4433 11203 4491 11209
rect 4433 11169 4445 11203
rect 4479 11169 4491 11203
rect 4433 11163 4491 11169
rect 4893 11203 4951 11209
rect 4893 11169 4905 11203
rect 4939 11200 4951 11203
rect 5074 11200 5080 11212
rect 4939 11172 5080 11200
rect 4939 11169 4951 11172
rect 4893 11163 4951 11169
rect 5074 11160 5080 11172
rect 5132 11160 5138 11212
rect 5166 11160 5172 11212
rect 5224 11200 5230 11212
rect 5442 11200 5448 11212
rect 5224 11172 5269 11200
rect 5403 11172 5448 11200
rect 5224 11160 5230 11172
rect 5442 11160 5448 11172
rect 5500 11160 5506 11212
rect 5994 11200 6000 11212
rect 5955 11172 6000 11200
rect 5994 11160 6000 11172
rect 6052 11160 6058 11212
rect 6454 11200 6460 11212
rect 6415 11172 6460 11200
rect 6454 11160 6460 11172
rect 6512 11160 6518 11212
rect 6730 11200 6736 11212
rect 6691 11172 6736 11200
rect 6730 11160 6736 11172
rect 6788 11160 6794 11212
rect 7006 11200 7012 11212
rect 6967 11172 7012 11200
rect 7006 11160 7012 11172
rect 7064 11160 7070 11212
rect 7190 11200 7196 11212
rect 7151 11172 7196 11200
rect 7190 11160 7196 11172
rect 7248 11160 7254 11212
rect 7926 11160 7932 11212
rect 7984 11200 7990 11212
rect 7984 11172 8248 11200
rect 7984 11160 7990 11172
rect 2958 11132 2964 11144
rect 2919 11104 2964 11132
rect 2958 11092 2964 11104
rect 3016 11092 3022 11144
rect 5261 11135 5319 11141
rect 5261 11101 5273 11135
rect 5307 11132 5319 11135
rect 6086 11132 6092 11144
rect 5307 11104 6092 11132
rect 5307 11101 5319 11104
rect 5261 11095 5319 11101
rect 6086 11092 6092 11104
rect 6144 11092 6150 11144
rect 6914 11132 6920 11144
rect 6875 11104 6920 11132
rect 6914 11092 6920 11104
rect 6972 11092 6978 11144
rect 8220 11141 8248 11172
rect 8662 11160 8668 11212
rect 8720 11200 8726 11212
rect 9861 11203 9919 11209
rect 9861 11200 9873 11203
rect 8720 11172 9873 11200
rect 8720 11160 8726 11172
rect 9861 11169 9873 11172
rect 9907 11169 9919 11203
rect 9861 11163 9919 11169
rect 9950 11160 9956 11212
rect 10008 11200 10014 11212
rect 10321 11203 10379 11209
rect 10008 11172 10053 11200
rect 10008 11160 10014 11172
rect 10321 11169 10333 11203
rect 10367 11200 10379 11203
rect 10778 11200 10784 11212
rect 10367 11172 10784 11200
rect 10367 11169 10379 11172
rect 10321 11163 10379 11169
rect 8205 11135 8263 11141
rect 8205 11101 8217 11135
rect 8251 11101 8263 11135
rect 8205 11095 8263 11101
rect 8846 11092 8852 11144
rect 8904 11132 8910 11144
rect 10336 11132 10364 11163
rect 10778 11160 10784 11172
rect 10836 11160 10842 11212
rect 11793 11203 11851 11209
rect 11793 11169 11805 11203
rect 11839 11200 11851 11203
rect 11974 11200 11980 11212
rect 11839 11172 11980 11200
rect 11839 11169 11851 11172
rect 11793 11163 11851 11169
rect 11974 11160 11980 11172
rect 12032 11160 12038 11212
rect 13262 11200 13268 11212
rect 13223 11172 13268 11200
rect 13262 11160 13268 11172
rect 13320 11160 13326 11212
rect 10594 11132 10600 11144
rect 8904 11104 10364 11132
rect 10428 11104 10600 11132
rect 8904 11092 8910 11104
rect 2406 11024 2412 11076
rect 2464 11064 2470 11076
rect 3053 11067 3111 11073
rect 3053 11064 3065 11067
rect 2464 11036 3065 11064
rect 2464 11024 2470 11036
rect 3053 11033 3065 11036
rect 3099 11033 3111 11067
rect 3053 11027 3111 11033
rect 4709 11067 4767 11073
rect 4709 11033 4721 11067
rect 4755 11064 4767 11067
rect 4798 11064 4804 11076
rect 4755 11036 4804 11064
rect 4755 11033 4767 11036
rect 4709 11027 4767 11033
rect 4798 11024 4804 11036
rect 4856 11024 4862 11076
rect 5718 11024 5724 11076
rect 5776 11064 5782 11076
rect 6822 11064 6828 11076
rect 5776 11036 6828 11064
rect 5776 11024 5782 11036
rect 6822 11024 6828 11036
rect 6880 11024 6886 11076
rect 9122 11024 9128 11076
rect 9180 11064 9186 11076
rect 10428 11064 10456 11104
rect 10594 11092 10600 11104
rect 10652 11132 10658 11144
rect 11149 11135 11207 11141
rect 11149 11132 11161 11135
rect 10652 11104 11161 11132
rect 10652 11092 10658 11104
rect 11149 11101 11161 11104
rect 11195 11101 11207 11135
rect 11149 11095 11207 11101
rect 9180 11036 10456 11064
rect 9180 11024 9186 11036
rect 5810 10956 5816 11008
rect 5868 10996 5874 11008
rect 9214 10996 9220 11008
rect 5868 10968 9220 10996
rect 5868 10956 5874 10968
rect 9214 10956 9220 10968
rect 9272 10956 9278 11008
rect 9858 10956 9864 11008
rect 9916 10996 9922 11008
rect 10060 11005 10088 11036
rect 10045 10999 10103 11005
rect 10045 10996 10057 10999
rect 9916 10968 10057 10996
rect 9916 10956 9922 10968
rect 10045 10965 10057 10968
rect 10091 10965 10103 10999
rect 10045 10959 10103 10965
rect 10137 10999 10195 11005
rect 10137 10965 10149 10999
rect 10183 10996 10195 10999
rect 10410 10996 10416 11008
rect 10183 10968 10416 10996
rect 10183 10965 10195 10968
rect 10137 10959 10195 10965
rect 10410 10956 10416 10968
rect 10468 10956 10474 11008
rect 10594 10996 10600 11008
rect 10555 10968 10600 10996
rect 10594 10956 10600 10968
rect 10652 10956 10658 11008
rect 1104 10906 13892 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 12246 10906
rect 12298 10854 12310 10906
rect 12362 10854 12374 10906
rect 12426 10854 12438 10906
rect 12490 10854 13892 10906
rect 1104 10832 13892 10854
rect 2869 10795 2927 10801
rect 2869 10761 2881 10795
rect 2915 10792 2927 10795
rect 2958 10792 2964 10804
rect 2915 10764 2964 10792
rect 2915 10761 2927 10764
rect 2869 10755 2927 10761
rect 2958 10752 2964 10764
rect 3016 10752 3022 10804
rect 5994 10792 6000 10804
rect 5828 10764 6000 10792
rect 4614 10724 4620 10736
rect 4575 10696 4620 10724
rect 4614 10684 4620 10696
rect 4672 10684 4678 10736
rect 2406 10656 2412 10668
rect 1596 10628 2412 10656
rect 1596 10597 1624 10628
rect 2406 10616 2412 10628
rect 2464 10616 2470 10668
rect 5258 10616 5264 10668
rect 5316 10656 5322 10668
rect 5537 10659 5595 10665
rect 5537 10656 5549 10659
rect 5316 10628 5549 10656
rect 5316 10616 5322 10628
rect 5537 10625 5549 10628
rect 5583 10625 5595 10659
rect 5828 10656 5856 10764
rect 5994 10752 6000 10764
rect 6052 10792 6058 10804
rect 6822 10792 6828 10804
rect 6052 10764 6828 10792
rect 6052 10752 6058 10764
rect 6822 10752 6828 10764
rect 6880 10752 6886 10804
rect 7834 10752 7840 10804
rect 7892 10792 7898 10804
rect 8665 10795 8723 10801
rect 8665 10792 8677 10795
rect 7892 10764 8677 10792
rect 7892 10752 7898 10764
rect 8665 10761 8677 10764
rect 8711 10792 8723 10795
rect 9309 10795 9367 10801
rect 9309 10792 9321 10795
rect 8711 10764 9321 10792
rect 8711 10761 8723 10764
rect 8665 10755 8723 10761
rect 9309 10761 9321 10764
rect 9355 10761 9367 10795
rect 9309 10755 9367 10761
rect 9582 10752 9588 10804
rect 9640 10792 9646 10804
rect 9677 10795 9735 10801
rect 9677 10792 9689 10795
rect 9640 10764 9689 10792
rect 9640 10752 9646 10764
rect 9677 10761 9689 10764
rect 9723 10761 9735 10795
rect 9677 10755 9735 10761
rect 11146 10752 11152 10804
rect 11204 10792 11210 10804
rect 11793 10795 11851 10801
rect 11793 10792 11805 10795
rect 11204 10764 11805 10792
rect 11204 10752 11210 10764
rect 11793 10761 11805 10764
rect 11839 10761 11851 10795
rect 11793 10755 11851 10761
rect 5905 10727 5963 10733
rect 5905 10693 5917 10727
rect 5951 10724 5963 10727
rect 12618 10724 12624 10736
rect 5951 10696 12624 10724
rect 5951 10693 5963 10696
rect 5905 10687 5963 10693
rect 12618 10684 12624 10696
rect 12676 10684 12682 10736
rect 7006 10656 7012 10668
rect 5537 10619 5595 10625
rect 5644 10628 5856 10656
rect 6967 10628 7012 10656
rect 1581 10591 1639 10597
rect 1581 10557 1593 10591
rect 1627 10557 1639 10591
rect 1854 10588 1860 10600
rect 1815 10560 1860 10588
rect 1581 10551 1639 10557
rect 1854 10548 1860 10560
rect 1912 10548 1918 10600
rect 2317 10591 2375 10597
rect 2317 10557 2329 10591
rect 2363 10588 2375 10591
rect 2682 10588 2688 10600
rect 2363 10560 2544 10588
rect 2643 10560 2688 10588
rect 2363 10557 2375 10560
rect 2317 10551 2375 10557
rect 1489 10523 1547 10529
rect 1489 10489 1501 10523
rect 1535 10520 1547 10523
rect 2409 10523 2467 10529
rect 2409 10520 2421 10523
rect 1535 10492 2421 10520
rect 1535 10489 1547 10492
rect 1489 10483 1547 10489
rect 2409 10489 2421 10492
rect 2455 10489 2467 10523
rect 2516 10520 2544 10560
rect 2682 10548 2688 10560
rect 2740 10548 2746 10600
rect 2774 10548 2780 10600
rect 2832 10588 2838 10600
rect 3145 10591 3203 10597
rect 3145 10588 3157 10591
rect 2832 10560 3157 10588
rect 2832 10548 2838 10560
rect 3145 10557 3157 10560
rect 3191 10557 3203 10591
rect 3145 10551 3203 10557
rect 4157 10591 4215 10597
rect 4157 10557 4169 10591
rect 4203 10557 4215 10591
rect 5442 10588 5448 10600
rect 5403 10560 5448 10588
rect 4157 10551 4215 10557
rect 2958 10520 2964 10532
rect 2516 10492 2964 10520
rect 2409 10483 2467 10489
rect 2958 10480 2964 10492
rect 3016 10520 3022 10532
rect 4062 10520 4068 10532
rect 3016 10492 4068 10520
rect 3016 10480 3022 10492
rect 4062 10480 4068 10492
rect 4120 10520 4126 10532
rect 4172 10520 4200 10551
rect 5442 10548 5448 10560
rect 5500 10548 5506 10600
rect 5644 10597 5672 10628
rect 7006 10616 7012 10628
rect 7064 10656 7070 10668
rect 7466 10656 7472 10668
rect 7064 10628 7472 10656
rect 7064 10616 7070 10628
rect 7466 10616 7472 10628
rect 7524 10616 7530 10668
rect 7561 10659 7619 10665
rect 7561 10625 7573 10659
rect 7607 10656 7619 10659
rect 7607 10628 8892 10656
rect 7607 10625 7619 10628
rect 7561 10619 7619 10625
rect 8864 10600 8892 10628
rect 9950 10616 9956 10668
rect 10008 10656 10014 10668
rect 10008 10628 10180 10656
rect 10008 10616 10014 10628
rect 5629 10591 5687 10597
rect 5629 10557 5641 10591
rect 5675 10557 5687 10591
rect 5629 10551 5687 10557
rect 5721 10591 5779 10597
rect 5721 10557 5733 10591
rect 5767 10588 5779 10591
rect 5902 10588 5908 10600
rect 5767 10560 5908 10588
rect 5767 10557 5779 10560
rect 5721 10551 5779 10557
rect 4120 10492 4200 10520
rect 4120 10480 4126 10492
rect 5350 10480 5356 10532
rect 5408 10520 5414 10532
rect 5644 10520 5672 10551
rect 5902 10548 5908 10560
rect 5960 10588 5966 10600
rect 7101 10591 7159 10597
rect 7101 10588 7113 10591
rect 5960 10560 7113 10588
rect 5960 10548 5966 10560
rect 7101 10557 7113 10560
rect 7147 10557 7159 10591
rect 7101 10551 7159 10557
rect 5408 10492 5672 10520
rect 5408 10480 5414 10492
rect 6730 10480 6736 10532
rect 6788 10520 6794 10532
rect 6825 10523 6883 10529
rect 6825 10520 6837 10523
rect 6788 10492 6837 10520
rect 6788 10480 6794 10492
rect 6825 10489 6837 10492
rect 6871 10489 6883 10523
rect 7116 10520 7144 10551
rect 7282 10548 7288 10600
rect 7340 10588 7346 10600
rect 7653 10591 7711 10597
rect 7653 10588 7665 10591
rect 7340 10560 7665 10588
rect 7340 10548 7346 10560
rect 7653 10557 7665 10560
rect 7699 10557 7711 10591
rect 7653 10551 7711 10557
rect 8665 10591 8723 10597
rect 8665 10557 8677 10591
rect 8711 10557 8723 10591
rect 8846 10588 8852 10600
rect 8807 10560 8852 10588
rect 8665 10551 8723 10557
rect 7561 10523 7619 10529
rect 7561 10520 7573 10523
rect 7116 10492 7573 10520
rect 6825 10483 6883 10489
rect 7561 10489 7573 10492
rect 7607 10489 7619 10523
rect 7834 10520 7840 10532
rect 7795 10492 7840 10520
rect 7561 10483 7619 10489
rect 7834 10480 7840 10492
rect 7892 10480 7898 10532
rect 7926 10480 7932 10532
rect 7984 10520 7990 10532
rect 8021 10523 8079 10529
rect 8021 10520 8033 10523
rect 7984 10492 8033 10520
rect 7984 10480 7990 10492
rect 8021 10489 8033 10492
rect 8067 10520 8079 10523
rect 8680 10520 8708 10551
rect 8846 10548 8852 10560
rect 8904 10548 8910 10600
rect 9306 10588 9312 10600
rect 9219 10560 9312 10588
rect 9306 10548 9312 10560
rect 9364 10588 9370 10600
rect 9401 10591 9459 10597
rect 9401 10588 9413 10591
rect 9364 10560 9413 10588
rect 9364 10548 9370 10560
rect 9401 10557 9413 10560
rect 9447 10557 9459 10591
rect 9401 10551 9459 10557
rect 9858 10548 9864 10600
rect 9916 10588 9922 10600
rect 10045 10591 10103 10597
rect 10045 10588 10057 10591
rect 9916 10560 10057 10588
rect 9916 10548 9922 10560
rect 10045 10557 10057 10560
rect 10091 10557 10103 10591
rect 10152 10588 10180 10628
rect 10226 10616 10232 10668
rect 10284 10656 10290 10668
rect 10502 10656 10508 10668
rect 10284 10628 10508 10656
rect 10284 10616 10290 10628
rect 10502 10616 10508 10628
rect 10560 10616 10566 10668
rect 10594 10616 10600 10668
rect 10652 10656 10658 10668
rect 10873 10659 10931 10665
rect 10873 10656 10885 10659
rect 10652 10628 10885 10656
rect 10652 10616 10658 10628
rect 10873 10625 10885 10628
rect 10919 10625 10931 10659
rect 10873 10619 10931 10625
rect 10962 10616 10968 10668
rect 11020 10656 11026 10668
rect 11020 10628 11744 10656
rect 11020 10616 11026 10628
rect 10413 10591 10471 10597
rect 10413 10588 10425 10591
rect 10152 10560 10425 10588
rect 10045 10551 10103 10557
rect 10413 10557 10425 10560
rect 10459 10557 10471 10591
rect 10413 10551 10471 10557
rect 11057 10591 11115 10597
rect 11057 10557 11069 10591
rect 11103 10588 11115 10591
rect 11146 10588 11152 10600
rect 11103 10560 11152 10588
rect 11103 10557 11115 10560
rect 11057 10551 11115 10557
rect 11146 10548 11152 10560
rect 11204 10548 11210 10600
rect 11716 10597 11744 10628
rect 11701 10591 11759 10597
rect 11701 10557 11713 10591
rect 11747 10557 11759 10591
rect 11701 10551 11759 10557
rect 11790 10548 11796 10600
rect 11848 10588 11854 10600
rect 11885 10591 11943 10597
rect 11885 10588 11897 10591
rect 11848 10560 11897 10588
rect 11848 10548 11854 10560
rect 11885 10557 11897 10560
rect 11931 10557 11943 10591
rect 12342 10588 12348 10600
rect 12303 10560 12348 10588
rect 11885 10551 11943 10557
rect 12342 10548 12348 10560
rect 12400 10548 12406 10600
rect 12986 10588 12992 10600
rect 12947 10560 12992 10588
rect 12986 10548 12992 10560
rect 13044 10548 13050 10600
rect 13262 10588 13268 10600
rect 13223 10560 13268 10588
rect 13262 10548 13268 10560
rect 13320 10548 13326 10600
rect 8067 10492 8708 10520
rect 8067 10489 8079 10492
rect 8021 10483 8079 10489
rect 9214 10480 9220 10532
rect 9272 10520 9278 10532
rect 9585 10523 9643 10529
rect 9585 10520 9597 10523
rect 9272 10492 9597 10520
rect 9272 10480 9278 10492
rect 9585 10489 9597 10492
rect 9631 10520 9643 10523
rect 10597 10523 10655 10529
rect 9631 10492 10548 10520
rect 9631 10489 9643 10492
rect 9585 10483 9643 10489
rect 3970 10412 3976 10464
rect 4028 10452 4034 10464
rect 7098 10452 7104 10464
rect 4028 10424 7104 10452
rect 4028 10412 4034 10424
rect 7098 10412 7104 10424
rect 7156 10412 7162 10464
rect 7285 10455 7343 10461
rect 7285 10421 7297 10455
rect 7331 10452 7343 10455
rect 7742 10452 7748 10464
rect 7331 10424 7748 10452
rect 7331 10421 7343 10424
rect 7285 10415 7343 10421
rect 7742 10412 7748 10424
rect 7800 10412 7806 10464
rect 9033 10455 9091 10461
rect 9033 10421 9045 10455
rect 9079 10452 9091 10455
rect 9950 10452 9956 10464
rect 9079 10424 9956 10452
rect 9079 10421 9091 10424
rect 9033 10415 9091 10421
rect 9950 10412 9956 10424
rect 10008 10412 10014 10464
rect 10244 10461 10272 10492
rect 10229 10455 10287 10461
rect 10229 10421 10241 10455
rect 10275 10421 10287 10455
rect 10229 10415 10287 10421
rect 10321 10455 10379 10461
rect 10321 10421 10333 10455
rect 10367 10452 10379 10455
rect 10410 10452 10416 10464
rect 10367 10424 10416 10452
rect 10367 10421 10379 10424
rect 10321 10415 10379 10421
rect 10410 10412 10416 10424
rect 10468 10412 10474 10464
rect 10520 10452 10548 10492
rect 10597 10489 10609 10523
rect 10643 10520 10655 10523
rect 11422 10520 11428 10532
rect 10643 10492 11428 10520
rect 10643 10489 10655 10492
rect 10597 10483 10655 10489
rect 11422 10480 11428 10492
rect 11480 10480 11486 10532
rect 11146 10452 11152 10464
rect 10520 10424 11152 10452
rect 11146 10412 11152 10424
rect 11204 10412 11210 10464
rect 11241 10455 11299 10461
rect 11241 10421 11253 10455
rect 11287 10452 11299 10455
rect 12526 10452 12532 10464
rect 11287 10424 12532 10452
rect 11287 10421 11299 10424
rect 11241 10415 11299 10421
rect 12526 10412 12532 10424
rect 12584 10412 12590 10464
rect 1104 10362 13892 10384
rect 1104 10310 8246 10362
rect 8298 10310 8310 10362
rect 8362 10310 8374 10362
rect 8426 10310 8438 10362
rect 8490 10310 13892 10362
rect 1104 10288 13892 10310
rect 5166 10208 5172 10260
rect 5224 10248 5230 10260
rect 5442 10248 5448 10260
rect 5224 10220 5448 10248
rect 5224 10208 5230 10220
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 6730 10248 6736 10260
rect 6643 10220 6736 10248
rect 2958 10180 2964 10192
rect 2919 10152 2964 10180
rect 2958 10140 2964 10152
rect 3016 10140 3022 10192
rect 4614 10180 4620 10192
rect 3344 10152 4620 10180
rect 1394 10112 1400 10124
rect 1307 10084 1400 10112
rect 1394 10072 1400 10084
rect 1452 10112 1458 10124
rect 1854 10112 1860 10124
rect 1452 10084 1860 10112
rect 1452 10072 1458 10084
rect 1854 10072 1860 10084
rect 1912 10072 1918 10124
rect 2682 10112 2688 10124
rect 2643 10084 2688 10112
rect 2682 10072 2688 10084
rect 2740 10072 2746 10124
rect 3344 10121 3372 10152
rect 4614 10140 4620 10152
rect 4672 10180 4678 10192
rect 4982 10180 4988 10192
rect 4672 10152 4988 10180
rect 4672 10140 4678 10152
rect 4982 10140 4988 10152
rect 5040 10140 5046 10192
rect 5810 10180 5816 10192
rect 5184 10152 5816 10180
rect 5184 10124 5212 10152
rect 5810 10140 5816 10152
rect 5868 10140 5874 10192
rect 3329 10115 3387 10121
rect 3329 10081 3341 10115
rect 3375 10081 3387 10115
rect 3329 10075 3387 10081
rect 3418 10072 3424 10124
rect 3476 10112 3482 10124
rect 3973 10115 4031 10121
rect 3973 10112 3985 10115
rect 3476 10084 3985 10112
rect 3476 10072 3482 10084
rect 3973 10081 3985 10084
rect 4019 10081 4031 10115
rect 3973 10075 4031 10081
rect 4249 10115 4307 10121
rect 4249 10081 4261 10115
rect 4295 10112 4307 10115
rect 4890 10112 4896 10124
rect 4295 10084 4896 10112
rect 4295 10081 4307 10084
rect 4249 10075 4307 10081
rect 4890 10072 4896 10084
rect 4948 10072 4954 10124
rect 5166 10112 5172 10124
rect 5079 10084 5172 10112
rect 5166 10072 5172 10084
rect 5224 10072 5230 10124
rect 5350 10072 5356 10124
rect 5408 10112 5414 10124
rect 5445 10115 5503 10121
rect 5445 10112 5457 10115
rect 5408 10084 5457 10112
rect 5408 10072 5414 10084
rect 5445 10081 5457 10084
rect 5491 10081 5503 10115
rect 5445 10075 5503 10081
rect 5537 10115 5595 10121
rect 5537 10081 5549 10115
rect 5583 10112 5595 10115
rect 5902 10112 5908 10124
rect 5583 10084 5908 10112
rect 5583 10081 5595 10084
rect 5537 10075 5595 10081
rect 5902 10072 5908 10084
rect 5960 10072 5966 10124
rect 6546 10112 6552 10124
rect 6507 10084 6552 10112
rect 6546 10072 6552 10084
rect 6604 10072 6610 10124
rect 6656 10112 6684 10220
rect 6730 10208 6736 10220
rect 6788 10248 6794 10260
rect 8754 10248 8760 10260
rect 6788 10220 8760 10248
rect 6788 10208 6794 10220
rect 6733 10115 6791 10121
rect 6733 10112 6745 10115
rect 6656 10084 6745 10112
rect 6733 10081 6745 10084
rect 6779 10081 6791 10115
rect 6914 10112 6920 10124
rect 6875 10084 6920 10112
rect 6733 10075 6791 10081
rect 6914 10072 6920 10084
rect 6972 10112 6978 10124
rect 7561 10115 7619 10121
rect 6972 10084 7512 10112
rect 6972 10072 6978 10084
rect 5261 10047 5319 10053
rect 5261 10013 5273 10047
rect 5307 10044 5319 10047
rect 5626 10044 5632 10056
rect 5307 10016 5632 10044
rect 5307 10013 5319 10016
rect 5261 10007 5319 10013
rect 5626 10004 5632 10016
rect 5684 10044 5690 10056
rect 6362 10044 6368 10056
rect 5684 10016 6368 10044
rect 5684 10004 5690 10016
rect 6362 10004 6368 10016
rect 6420 10004 6426 10056
rect 6638 10004 6644 10056
rect 6696 10044 6702 10056
rect 7377 10047 7435 10053
rect 7377 10044 7389 10047
rect 6696 10016 7389 10044
rect 6696 10004 6702 10016
rect 7377 10013 7389 10016
rect 7423 10013 7435 10047
rect 7484 10044 7512 10084
rect 7561 10081 7573 10115
rect 7607 10112 7619 10115
rect 7668 10112 7696 10220
rect 8754 10208 8760 10220
rect 8812 10248 8818 10260
rect 10045 10251 10103 10257
rect 10045 10248 10057 10251
rect 8812 10220 10057 10248
rect 8812 10208 8818 10220
rect 10045 10217 10057 10220
rect 10091 10248 10103 10251
rect 10134 10248 10140 10260
rect 10091 10220 10140 10248
rect 10091 10217 10103 10220
rect 10045 10211 10103 10217
rect 10134 10208 10140 10220
rect 10192 10248 10198 10260
rect 11698 10248 11704 10260
rect 10192 10220 11704 10248
rect 10192 10208 10198 10220
rect 11698 10208 11704 10220
rect 11756 10208 11762 10260
rect 9217 10183 9275 10189
rect 9217 10149 9229 10183
rect 9263 10180 9275 10183
rect 10226 10180 10232 10192
rect 9263 10152 10232 10180
rect 9263 10149 9275 10152
rect 9217 10143 9275 10149
rect 10226 10140 10232 10152
rect 10284 10140 10290 10192
rect 10594 10180 10600 10192
rect 10428 10152 10600 10180
rect 7607 10084 7696 10112
rect 7607 10081 7619 10084
rect 7561 10075 7619 10081
rect 7742 10072 7748 10124
rect 7800 10112 7806 10124
rect 7837 10115 7895 10121
rect 7837 10112 7849 10115
rect 7800 10084 7849 10112
rect 7800 10072 7806 10084
rect 7837 10081 7849 10084
rect 7883 10081 7895 10115
rect 8018 10112 8024 10124
rect 7979 10084 8024 10112
rect 7837 10075 7895 10081
rect 8018 10072 8024 10084
rect 8076 10072 8082 10124
rect 8110 10072 8116 10124
rect 8168 10112 8174 10124
rect 8297 10115 8355 10121
rect 8297 10112 8309 10115
rect 8168 10084 8309 10112
rect 8168 10072 8174 10084
rect 8297 10081 8309 10084
rect 8343 10081 8355 10115
rect 8570 10112 8576 10124
rect 8531 10084 8576 10112
rect 8297 10075 8355 10081
rect 8570 10072 8576 10084
rect 8628 10072 8634 10124
rect 8662 10072 8668 10124
rect 8720 10112 8726 10124
rect 9125 10115 9183 10121
rect 9125 10112 9137 10115
rect 8720 10084 9137 10112
rect 8720 10072 8726 10084
rect 9125 10081 9137 10084
rect 9171 10081 9183 10115
rect 9306 10112 9312 10124
rect 9267 10084 9312 10112
rect 9125 10075 9183 10081
rect 9306 10072 9312 10084
rect 9364 10072 9370 10124
rect 9490 10112 9496 10124
rect 9451 10084 9496 10112
rect 9490 10072 9496 10084
rect 9548 10072 9554 10124
rect 9766 10072 9772 10124
rect 9824 10112 9830 10124
rect 10428 10121 10456 10152
rect 10594 10140 10600 10152
rect 10652 10140 10658 10192
rect 12710 10180 12716 10192
rect 11914 10152 12716 10180
rect 12710 10140 12716 10152
rect 12768 10140 12774 10192
rect 13078 10180 13084 10192
rect 13039 10152 13084 10180
rect 13078 10140 13084 10152
rect 13136 10140 13142 10192
rect 9953 10115 10011 10121
rect 9953 10112 9965 10115
rect 9824 10084 9965 10112
rect 9824 10072 9830 10084
rect 9953 10081 9965 10084
rect 9999 10081 10011 10115
rect 9953 10075 10011 10081
rect 10413 10115 10471 10121
rect 10413 10081 10425 10115
rect 10459 10081 10471 10115
rect 12986 10112 12992 10124
rect 12947 10084 12992 10112
rect 10413 10075 10471 10081
rect 12986 10072 12992 10084
rect 13044 10072 13050 10124
rect 8588 10044 8616 10072
rect 8754 10044 8760 10056
rect 7484 10016 7788 10044
rect 8588 10016 8760 10044
rect 7377 10007 7435 10013
rect 3970 9976 3976 9988
rect 3931 9948 3976 9976
rect 3970 9936 3976 9948
rect 4028 9936 4034 9988
rect 4062 9936 4068 9988
rect 4120 9976 4126 9988
rect 7760 9985 7788 10016
rect 8754 10004 8760 10016
rect 8812 10004 8818 10056
rect 10686 10044 10692 10056
rect 10647 10016 10692 10044
rect 10686 10004 10692 10016
rect 10744 10004 10750 10056
rect 12066 10004 12072 10056
rect 12124 10044 12130 10056
rect 12342 10044 12348 10056
rect 12124 10016 12348 10044
rect 12124 10004 12130 10016
rect 12342 10004 12348 10016
rect 12400 10044 12406 10056
rect 12529 10047 12587 10053
rect 12529 10044 12541 10047
rect 12400 10016 12541 10044
rect 12400 10004 12406 10016
rect 12529 10013 12541 10016
rect 12575 10013 12587 10047
rect 12529 10007 12587 10013
rect 6273 9979 6331 9985
rect 6273 9976 6285 9979
rect 4120 9948 6285 9976
rect 4120 9936 4126 9948
rect 6273 9945 6285 9948
rect 6319 9945 6331 9979
rect 7653 9979 7711 9985
rect 7653 9976 7665 9979
rect 6273 9939 6331 9945
rect 6656 9948 7665 9976
rect 3513 9911 3571 9917
rect 3513 9877 3525 9911
rect 3559 9908 3571 9911
rect 4614 9908 4620 9920
rect 3559 9880 4620 9908
rect 3559 9877 3571 9880
rect 3513 9871 3571 9877
rect 4614 9868 4620 9880
rect 4672 9868 4678 9920
rect 4890 9908 4896 9920
rect 4851 9880 4896 9908
rect 4890 9868 4896 9880
rect 4948 9868 4954 9920
rect 5353 9911 5411 9917
rect 5353 9877 5365 9911
rect 5399 9908 5411 9911
rect 5442 9908 5448 9920
rect 5399 9880 5448 9908
rect 5399 9877 5411 9880
rect 5353 9871 5411 9877
rect 5442 9868 5448 9880
rect 5500 9868 5506 9920
rect 5810 9868 5816 9920
rect 5868 9908 5874 9920
rect 6086 9908 6092 9920
rect 5868 9880 6092 9908
rect 5868 9868 5874 9880
rect 6086 9868 6092 9880
rect 6144 9908 6150 9920
rect 6656 9917 6684 9948
rect 7653 9945 7665 9948
rect 7699 9945 7711 9979
rect 7653 9939 7711 9945
rect 7745 9979 7803 9985
rect 7745 9945 7757 9979
rect 7791 9976 7803 9979
rect 7834 9976 7840 9988
rect 7791 9948 7840 9976
rect 7791 9945 7803 9948
rect 7745 9939 7803 9945
rect 7834 9936 7840 9948
rect 7892 9936 7898 9988
rect 8570 9976 8576 9988
rect 8531 9948 8576 9976
rect 8570 9936 8576 9948
rect 8628 9936 8634 9988
rect 6641 9911 6699 9917
rect 6641 9908 6653 9911
rect 6144 9880 6653 9908
rect 6144 9868 6150 9880
rect 6641 9877 6653 9880
rect 6687 9877 6699 9911
rect 6641 9871 6699 9877
rect 6825 9911 6883 9917
rect 6825 9877 6837 9911
rect 6871 9908 6883 9911
rect 7374 9908 7380 9920
rect 6871 9880 7380 9908
rect 6871 9877 6883 9880
rect 6825 9871 6883 9877
rect 7374 9868 7380 9880
rect 7432 9868 7438 9920
rect 11974 9868 11980 9920
rect 12032 9908 12038 9920
rect 12161 9911 12219 9917
rect 12161 9908 12173 9911
rect 12032 9880 12173 9908
rect 12032 9868 12038 9880
rect 12161 9877 12173 9880
rect 12207 9877 12219 9911
rect 12161 9871 12219 9877
rect 1104 9818 13892 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 12246 9818
rect 12298 9766 12310 9818
rect 12362 9766 12374 9818
rect 12426 9766 12438 9818
rect 12490 9766 13892 9818
rect 1104 9744 13892 9766
rect 1394 9704 1400 9716
rect 1355 9676 1400 9704
rect 1394 9664 1400 9676
rect 1452 9664 1458 9716
rect 3326 9704 3332 9716
rect 3287 9676 3332 9704
rect 3326 9664 3332 9676
rect 3384 9664 3390 9716
rect 5534 9704 5540 9716
rect 5495 9676 5540 9704
rect 5534 9664 5540 9676
rect 5592 9664 5598 9716
rect 5718 9704 5724 9716
rect 5679 9676 5724 9704
rect 5718 9664 5724 9676
rect 5776 9664 5782 9716
rect 7006 9664 7012 9716
rect 7064 9704 7070 9716
rect 7101 9707 7159 9713
rect 7101 9704 7113 9707
rect 7064 9676 7113 9704
rect 7064 9664 7070 9676
rect 7101 9673 7113 9676
rect 7147 9673 7159 9707
rect 9214 9704 9220 9716
rect 7101 9667 7159 9673
rect 8266 9676 9220 9704
rect 4890 9636 4896 9648
rect 1780 9608 4896 9636
rect 1780 9509 1808 9608
rect 4890 9596 4896 9608
rect 4948 9596 4954 9648
rect 6822 9596 6828 9648
rect 6880 9636 6886 9648
rect 8266 9636 8294 9676
rect 9214 9664 9220 9676
rect 9272 9704 9278 9716
rect 10410 9704 10416 9716
rect 9272 9676 10416 9704
rect 9272 9664 9278 9676
rect 10410 9664 10416 9676
rect 10468 9664 10474 9716
rect 10686 9664 10692 9716
rect 10744 9704 10750 9716
rect 10781 9707 10839 9713
rect 10781 9704 10793 9707
rect 10744 9676 10793 9704
rect 10744 9664 10750 9676
rect 10781 9673 10793 9676
rect 10827 9673 10839 9707
rect 10781 9667 10839 9673
rect 12066 9664 12072 9716
rect 12124 9704 12130 9716
rect 12253 9707 12311 9713
rect 12253 9704 12265 9707
rect 12124 9676 12265 9704
rect 12124 9664 12130 9676
rect 12253 9673 12265 9676
rect 12299 9673 12311 9707
rect 12253 9667 12311 9673
rect 8938 9636 8944 9648
rect 6880 9608 8294 9636
rect 8899 9608 8944 9636
rect 6880 9596 6886 9608
rect 2038 9568 2044 9580
rect 1999 9540 2044 9568
rect 2038 9528 2044 9540
rect 2096 9528 2102 9580
rect 5626 9528 5632 9580
rect 5684 9568 5690 9580
rect 8266 9577 8294 9608
rect 8938 9596 8944 9608
rect 8996 9596 9002 9648
rect 9122 9636 9128 9648
rect 9048 9608 9128 9636
rect 6641 9571 6699 9577
rect 6641 9568 6653 9571
rect 5684 9540 6653 9568
rect 5684 9528 5690 9540
rect 6641 9537 6653 9540
rect 6687 9537 6699 9571
rect 8266 9571 8335 9577
rect 8266 9540 8289 9571
rect 6641 9531 6699 9537
rect 8277 9537 8289 9540
rect 8323 9537 8335 9571
rect 8277 9531 8335 9537
rect 1765 9503 1823 9509
rect 1765 9469 1777 9503
rect 1811 9469 1823 9503
rect 1765 9463 1823 9469
rect 2777 9503 2835 9509
rect 2777 9469 2789 9503
rect 2823 9500 2835 9503
rect 2866 9500 2872 9512
rect 2823 9472 2872 9500
rect 2823 9469 2835 9472
rect 2777 9463 2835 9469
rect 2866 9460 2872 9472
rect 2924 9460 2930 9512
rect 3234 9500 3240 9512
rect 3195 9472 3240 9500
rect 3234 9460 3240 9472
rect 3292 9460 3298 9512
rect 3510 9500 3516 9512
rect 3471 9472 3516 9500
rect 3510 9460 3516 9472
rect 3568 9460 3574 9512
rect 4614 9500 4620 9512
rect 4575 9472 4620 9500
rect 4614 9460 4620 9472
rect 4672 9460 4678 9512
rect 5258 9460 5264 9512
rect 5316 9500 5322 9512
rect 6733 9503 6791 9509
rect 5316 9472 6040 9500
rect 5316 9460 5322 9472
rect 3602 9392 3608 9444
rect 3660 9432 3666 9444
rect 3973 9435 4031 9441
rect 3973 9432 3985 9435
rect 3660 9404 3985 9432
rect 3660 9392 3666 9404
rect 3973 9401 3985 9404
rect 4019 9432 4031 9435
rect 5626 9432 5632 9444
rect 4019 9404 5632 9432
rect 4019 9401 4031 9404
rect 3973 9395 4031 9401
rect 5626 9392 5632 9404
rect 5684 9392 5690 9444
rect 5721 9435 5779 9441
rect 5721 9401 5733 9435
rect 5767 9432 5779 9435
rect 5810 9432 5816 9444
rect 5767 9404 5816 9432
rect 5767 9401 5779 9404
rect 5721 9395 5779 9401
rect 5810 9392 5816 9404
rect 5868 9392 5874 9444
rect 5905 9435 5963 9441
rect 5905 9401 5917 9435
rect 5951 9401 5963 9435
rect 6012 9432 6040 9472
rect 6733 9469 6745 9503
rect 6779 9500 6791 9503
rect 7926 9500 7932 9512
rect 6779 9472 7932 9500
rect 6779 9469 6791 9472
rect 6733 9463 6791 9469
rect 7926 9460 7932 9472
rect 7984 9460 7990 9512
rect 9048 9509 9076 9608
rect 9122 9596 9128 9608
rect 9180 9636 9186 9648
rect 9861 9639 9919 9645
rect 9861 9636 9873 9639
rect 9180 9608 9873 9636
rect 9180 9596 9186 9608
rect 9861 9605 9873 9608
rect 9907 9605 9919 9639
rect 9861 9599 9919 9605
rect 9769 9571 9827 9577
rect 9769 9537 9781 9571
rect 9815 9568 9827 9571
rect 10778 9568 10784 9580
rect 9815 9540 10784 9568
rect 9815 9537 9827 9540
rect 9769 9531 9827 9537
rect 10778 9528 10784 9540
rect 10836 9568 10842 9580
rect 11241 9571 11299 9577
rect 11241 9568 11253 9571
rect 10836 9540 11253 9568
rect 10836 9528 10842 9540
rect 11241 9537 11253 9540
rect 11287 9568 11299 9571
rect 11793 9571 11851 9577
rect 11793 9568 11805 9571
rect 11287 9540 11805 9568
rect 11287 9537 11299 9540
rect 11241 9531 11299 9537
rect 11793 9537 11805 9540
rect 11839 9537 11851 9571
rect 12802 9568 12808 9580
rect 12763 9540 12808 9568
rect 11793 9531 11851 9537
rect 12802 9528 12808 9540
rect 12860 9528 12866 9580
rect 8573 9503 8631 9509
rect 8573 9469 8585 9503
rect 8619 9500 8631 9503
rect 9048 9503 9131 9509
rect 8619 9472 8984 9500
rect 9048 9472 9085 9503
rect 8619 9469 8631 9472
rect 8573 9463 8631 9469
rect 7193 9435 7251 9441
rect 7193 9432 7205 9435
rect 6012 9404 7205 9432
rect 5905 9395 5963 9401
rect 7193 9401 7205 9404
rect 7239 9401 7251 9435
rect 7374 9432 7380 9444
rect 7335 9404 7380 9432
rect 7193 9395 7251 9401
rect 1486 9324 1492 9376
rect 1544 9364 1550 9376
rect 1857 9367 1915 9373
rect 1857 9364 1869 9367
rect 1544 9336 1869 9364
rect 1544 9324 1550 9336
rect 1857 9333 1869 9336
rect 1903 9333 1915 9367
rect 1857 9327 1915 9333
rect 2774 9324 2780 9376
rect 2832 9364 2838 9376
rect 2869 9367 2927 9373
rect 2869 9364 2881 9367
rect 2832 9336 2881 9364
rect 2832 9324 2838 9336
rect 2869 9333 2881 9336
rect 2915 9333 2927 9367
rect 2869 9327 2927 9333
rect 5442 9324 5448 9376
rect 5500 9364 5506 9376
rect 5920 9364 5948 9395
rect 7374 9392 7380 9404
rect 7432 9392 7438 9444
rect 7466 9392 7472 9444
rect 7524 9432 7530 9444
rect 7837 9435 7895 9441
rect 7837 9432 7849 9435
rect 7524 9404 7849 9432
rect 7524 9392 7530 9404
rect 7837 9401 7849 9404
rect 7883 9401 7895 9435
rect 7837 9395 7895 9401
rect 8021 9435 8079 9441
rect 8021 9401 8033 9435
rect 8067 9432 8079 9435
rect 8110 9432 8116 9444
rect 8067 9404 8116 9432
rect 8067 9401 8079 9404
rect 8021 9395 8079 9401
rect 8110 9392 8116 9404
rect 8168 9392 8174 9444
rect 8481 9435 8539 9441
rect 8481 9401 8493 9435
rect 8527 9432 8539 9435
rect 8662 9432 8668 9444
rect 8527 9404 8668 9432
rect 8527 9401 8539 9404
rect 8481 9395 8539 9401
rect 8662 9392 8668 9404
rect 8720 9392 8726 9444
rect 7006 9364 7012 9376
rect 5500 9336 7012 9364
rect 5500 9324 5506 9336
rect 7006 9324 7012 9336
rect 7064 9324 7070 9376
rect 7926 9324 7932 9376
rect 7984 9364 7990 9376
rect 8389 9367 8447 9373
rect 8389 9364 8401 9367
rect 7984 9336 8401 9364
rect 7984 9324 7990 9336
rect 8389 9333 8401 9336
rect 8435 9333 8447 9367
rect 8956 9364 8984 9472
rect 9073 9469 9085 9472
rect 9119 9469 9131 9503
rect 9073 9463 9131 9469
rect 9214 9460 9220 9512
rect 9272 9500 9278 9512
rect 9490 9500 9496 9512
rect 9272 9472 9316 9500
rect 9451 9472 9496 9500
rect 9272 9460 9278 9472
rect 9490 9460 9496 9472
rect 9548 9460 9554 9512
rect 10045 9503 10103 9509
rect 10045 9469 10057 9503
rect 10091 9469 10103 9503
rect 10045 9463 10103 9469
rect 10137 9503 10195 9509
rect 10137 9469 10149 9503
rect 10183 9500 10195 9503
rect 10183 9472 10921 9500
rect 10183 9469 10195 9472
rect 10137 9463 10195 9469
rect 9306 9392 9312 9444
rect 9364 9432 9370 9444
rect 9508 9432 9536 9460
rect 10060 9432 10088 9463
rect 9364 9404 9409 9432
rect 9508 9404 10088 9432
rect 10689 9435 10747 9441
rect 9364 9392 9370 9404
rect 10689 9401 10701 9435
rect 10735 9401 10747 9435
rect 10893 9432 10921 9472
rect 10962 9460 10968 9512
rect 11020 9500 11026 9512
rect 11057 9503 11115 9509
rect 11057 9500 11069 9503
rect 11020 9472 11069 9500
rect 11020 9460 11026 9472
rect 11057 9469 11069 9472
rect 11103 9469 11115 9503
rect 11057 9463 11115 9469
rect 11885 9503 11943 9509
rect 11885 9469 11897 9503
rect 11931 9500 11943 9503
rect 11974 9500 11980 9512
rect 11931 9472 11980 9500
rect 11931 9469 11943 9472
rect 11885 9463 11943 9469
rect 11146 9432 11152 9444
rect 10893 9404 11152 9432
rect 10689 9395 10747 9401
rect 9858 9364 9864 9376
rect 8956 9336 9864 9364
rect 8389 9327 8447 9333
rect 9858 9324 9864 9336
rect 9916 9324 9922 9376
rect 10321 9367 10379 9373
rect 10321 9333 10333 9367
rect 10367 9364 10379 9367
rect 10410 9364 10416 9376
rect 10367 9336 10416 9364
rect 10367 9333 10379 9336
rect 10321 9327 10379 9333
rect 10410 9324 10416 9336
rect 10468 9324 10474 9376
rect 10704 9364 10732 9395
rect 11146 9392 11152 9404
rect 11204 9432 11210 9444
rect 11900 9432 11928 9463
rect 11974 9460 11980 9472
rect 12032 9460 12038 9512
rect 12618 9500 12624 9512
rect 12579 9472 12624 9500
rect 12618 9460 12624 9472
rect 12676 9460 12682 9512
rect 11204 9404 11928 9432
rect 11204 9392 11210 9404
rect 10778 9364 10784 9376
rect 10704 9336 10784 9364
rect 10778 9324 10784 9336
rect 10836 9324 10842 9376
rect 12713 9367 12771 9373
rect 12713 9333 12725 9367
rect 12759 9364 12771 9367
rect 13814 9364 13820 9376
rect 12759 9336 13820 9364
rect 12759 9333 12771 9336
rect 12713 9327 12771 9333
rect 13814 9324 13820 9336
rect 13872 9324 13878 9376
rect 1104 9274 13892 9296
rect 1104 9222 8246 9274
rect 8298 9222 8310 9274
rect 8362 9222 8374 9274
rect 8426 9222 8438 9274
rect 8490 9222 13892 9274
rect 1104 9200 13892 9222
rect 1949 9163 2007 9169
rect 1949 9129 1961 9163
rect 1995 9160 2007 9163
rect 2685 9163 2743 9169
rect 1995 9132 2636 9160
rect 1995 9129 2007 9132
rect 1949 9123 2007 9129
rect 1581 9095 1639 9101
rect 1581 9061 1593 9095
rect 1627 9092 1639 9095
rect 2608 9092 2636 9132
rect 2685 9129 2697 9163
rect 2731 9160 2743 9163
rect 4249 9163 4307 9169
rect 2731 9132 4200 9160
rect 2731 9129 2743 9132
rect 2685 9123 2743 9129
rect 3050 9092 3056 9104
rect 1627 9064 2544 9092
rect 2608 9064 3056 9092
rect 1627 9061 1639 9064
rect 1581 9055 1639 9061
rect 1857 9027 1915 9033
rect 1857 8993 1869 9027
rect 1903 9024 1915 9027
rect 2130 9024 2136 9036
rect 1903 8996 2136 9024
rect 1903 8993 1915 8996
rect 1857 8987 1915 8993
rect 2130 8984 2136 8996
rect 2188 8984 2194 9036
rect 2314 9024 2320 9036
rect 2275 8996 2320 9024
rect 2314 8984 2320 8996
rect 2372 8984 2378 9036
rect 2516 9024 2544 9064
rect 3050 9052 3056 9064
rect 3108 9052 3114 9104
rect 3326 9052 3332 9104
rect 3384 9092 3390 9104
rect 4172 9092 4200 9132
rect 4249 9129 4261 9163
rect 4295 9160 4307 9163
rect 4982 9160 4988 9172
rect 4295 9132 4988 9160
rect 4295 9129 4307 9132
rect 4249 9123 4307 9129
rect 4982 9120 4988 9132
rect 5040 9120 5046 9172
rect 5166 9120 5172 9172
rect 5224 9160 5230 9172
rect 5534 9160 5540 9172
rect 5224 9132 5540 9160
rect 5224 9120 5230 9132
rect 5534 9120 5540 9132
rect 5592 9160 5598 9172
rect 6822 9160 6828 9172
rect 5592 9132 6828 9160
rect 5592 9120 5598 9132
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 9490 9160 9496 9172
rect 7852 9132 9496 9160
rect 5258 9092 5264 9104
rect 3384 9064 3924 9092
rect 4172 9064 5264 9092
rect 3384 9052 3390 9064
rect 3896 9033 3924 9064
rect 5258 9052 5264 9064
rect 5316 9052 5322 9104
rect 6086 9052 6092 9104
rect 6144 9052 6150 9104
rect 7101 9095 7159 9101
rect 7101 9061 7113 9095
rect 7147 9092 7159 9095
rect 7466 9092 7472 9104
rect 7147 9064 7472 9092
rect 7147 9061 7159 9064
rect 7101 9055 7159 9061
rect 7466 9052 7472 9064
rect 7524 9052 7530 9104
rect 3881 9027 3939 9033
rect 2516 8996 3832 9024
rect 2685 8959 2743 8965
rect 2685 8956 2697 8959
rect 2424 8928 2697 8956
rect 1489 8891 1547 8897
rect 1489 8857 1501 8891
rect 1535 8888 1547 8891
rect 2424 8888 2452 8928
rect 2685 8925 2697 8928
rect 2731 8925 2743 8959
rect 2685 8919 2743 8925
rect 2777 8959 2835 8965
rect 2777 8925 2789 8959
rect 2823 8925 2835 8959
rect 3326 8956 3332 8968
rect 3287 8928 3332 8956
rect 2777 8919 2835 8925
rect 1535 8860 2452 8888
rect 2501 8891 2559 8897
rect 1535 8857 1547 8860
rect 1489 8851 1547 8857
rect 2501 8857 2513 8891
rect 2547 8888 2559 8891
rect 2792 8888 2820 8919
rect 3326 8916 3332 8928
rect 3384 8916 3390 8968
rect 3804 8956 3832 8996
rect 3881 8993 3893 9027
rect 3927 8993 3939 9027
rect 3881 8987 3939 8993
rect 4249 9027 4307 9033
rect 4249 8993 4261 9027
rect 4295 9024 4307 9027
rect 4706 9024 4712 9036
rect 4295 8996 4712 9024
rect 4295 8993 4307 8996
rect 4249 8987 4307 8993
rect 4706 8984 4712 8996
rect 4764 8984 4770 9036
rect 4890 9024 4896 9036
rect 4851 8996 4896 9024
rect 4890 8984 4896 8996
rect 4948 8984 4954 9036
rect 4985 9027 5043 9033
rect 4985 8993 4997 9027
rect 5031 8993 5043 9027
rect 5166 9024 5172 9036
rect 5127 8996 5172 9024
rect 4985 8987 5043 8993
rect 4614 8956 4620 8968
rect 3804 8928 4620 8956
rect 4614 8916 4620 8928
rect 4672 8916 4678 8968
rect 5000 8956 5028 8987
rect 5166 8984 5172 8996
rect 5224 8984 5230 9036
rect 7558 8984 7564 9036
rect 7616 9024 7622 9036
rect 7852 9033 7880 9132
rect 8754 9092 8760 9104
rect 8036 9064 8760 9092
rect 8036 9033 8064 9064
rect 8754 9052 8760 9064
rect 8812 9052 8818 9104
rect 9232 9036 9260 9132
rect 9490 9120 9496 9132
rect 9548 9120 9554 9172
rect 9582 9120 9588 9172
rect 9640 9160 9646 9172
rect 9953 9163 10011 9169
rect 9953 9160 9965 9163
rect 9640 9132 9965 9160
rect 9640 9120 9646 9132
rect 9953 9129 9965 9132
rect 9999 9129 10011 9163
rect 10778 9160 10784 9172
rect 10739 9132 10784 9160
rect 9953 9123 10011 9129
rect 10778 9120 10784 9132
rect 10836 9120 10842 9172
rect 11057 9163 11115 9169
rect 11057 9129 11069 9163
rect 11103 9160 11115 9163
rect 12710 9160 12716 9172
rect 11103 9132 12296 9160
rect 12671 9132 12716 9160
rect 11103 9129 11115 9132
rect 11057 9123 11115 9129
rect 9398 9092 9404 9104
rect 9324 9064 9404 9092
rect 7837 9027 7895 9033
rect 7837 9024 7849 9027
rect 7616 8996 7849 9024
rect 7616 8984 7622 8996
rect 7837 8993 7849 8996
rect 7883 8993 7895 9027
rect 7837 8987 7895 8993
rect 8021 9027 8079 9033
rect 8021 8993 8033 9027
rect 8067 8993 8079 9027
rect 8021 8987 8079 8993
rect 8297 9027 8355 9033
rect 8297 8993 8309 9027
rect 8343 9024 8355 9027
rect 8570 9024 8576 9036
rect 8343 8996 8576 9024
rect 8343 8993 8355 8996
rect 8297 8987 8355 8993
rect 8570 8984 8576 8996
rect 8628 8984 8634 9036
rect 9125 9027 9183 9033
rect 9125 8993 9137 9027
rect 9171 9024 9183 9027
rect 9214 9024 9220 9036
rect 9171 8996 9220 9024
rect 9171 8993 9183 8996
rect 9125 8987 9183 8993
rect 9214 8984 9220 8996
rect 9272 8984 9278 9036
rect 9324 9033 9352 9064
rect 9398 9052 9404 9064
rect 9456 9052 9462 9104
rect 10410 9092 10416 9104
rect 9646 9064 10416 9092
rect 9309 9027 9367 9033
rect 9309 8993 9321 9027
rect 9355 8993 9367 9027
rect 9309 8987 9367 8993
rect 9493 9027 9551 9033
rect 9493 8993 9505 9027
rect 9539 9024 9551 9027
rect 9646 9024 9674 9064
rect 10410 9052 10416 9064
rect 10468 9052 10474 9104
rect 10505 9095 10563 9101
rect 10505 9061 10517 9095
rect 10551 9092 10563 9095
rect 11885 9095 11943 9101
rect 11885 9092 11897 9095
rect 10551 9064 11897 9092
rect 10551 9061 10563 9064
rect 10505 9055 10563 9061
rect 11885 9061 11897 9064
rect 11931 9061 11943 9095
rect 11885 9055 11943 9061
rect 9539 8996 9674 9024
rect 9953 9027 10011 9033
rect 9539 8993 9551 8996
rect 9493 8987 9551 8993
rect 9953 8993 9965 9027
rect 9999 9024 10011 9027
rect 10137 9027 10195 9033
rect 10137 9024 10149 9027
rect 9999 8996 10149 9024
rect 9999 8993 10011 8996
rect 9953 8987 10011 8993
rect 10137 8993 10149 8996
rect 10183 8993 10195 9027
rect 10137 8987 10195 8993
rect 10285 9027 10343 9033
rect 10285 8993 10297 9027
rect 10331 8993 10343 9027
rect 10285 8987 10343 8993
rect 5629 8959 5687 8965
rect 5629 8956 5641 8959
rect 5000 8928 5641 8956
rect 5629 8925 5641 8928
rect 5675 8925 5687 8959
rect 7377 8959 7435 8965
rect 7377 8956 7389 8959
rect 5629 8919 5687 8925
rect 6104 8928 7389 8956
rect 2547 8860 2820 8888
rect 2547 8857 2559 8860
rect 2501 8851 2559 8857
rect 2866 8848 2872 8900
rect 2924 8888 2930 8900
rect 5077 8891 5135 8897
rect 2924 8860 2969 8888
rect 2924 8848 2930 8860
rect 5077 8857 5089 8891
rect 5123 8888 5135 8891
rect 5442 8888 5448 8900
rect 5123 8860 5448 8888
rect 5123 8857 5135 8860
rect 5077 8851 5135 8857
rect 5442 8848 5448 8860
rect 5500 8848 5506 8900
rect 1762 8780 1768 8832
rect 1820 8820 1826 8832
rect 4709 8823 4767 8829
rect 4709 8820 4721 8823
rect 1820 8792 4721 8820
rect 1820 8780 1826 8792
rect 4709 8789 4721 8792
rect 4755 8789 4767 8823
rect 5644 8820 5672 8919
rect 5718 8848 5724 8900
rect 5776 8888 5782 8900
rect 6104 8888 6132 8928
rect 7377 8925 7389 8928
rect 7423 8956 7435 8959
rect 7466 8956 7472 8968
rect 7423 8928 7472 8956
rect 7423 8925 7435 8928
rect 7377 8919 7435 8925
rect 7466 8916 7472 8928
rect 7524 8916 7530 8968
rect 8113 8959 8171 8965
rect 8113 8925 8125 8959
rect 8159 8925 8171 8959
rect 8113 8919 8171 8925
rect 5776 8860 6132 8888
rect 5776 8848 5782 8860
rect 7834 8848 7840 8900
rect 7892 8888 7898 8900
rect 8128 8888 8156 8919
rect 8202 8916 8208 8968
rect 8260 8956 8266 8968
rect 9401 8959 9459 8965
rect 9401 8956 9413 8959
rect 8260 8928 8305 8956
rect 8772 8928 9413 8956
rect 8260 8916 8266 8928
rect 8772 8900 8800 8928
rect 9401 8925 9413 8928
rect 9447 8925 9459 8959
rect 9401 8919 9459 8925
rect 9586 8959 9644 8965
rect 9586 8925 9598 8959
rect 9632 8925 9644 8959
rect 10300 8956 10328 8987
rect 10594 8984 10600 9036
rect 10652 9033 10658 9036
rect 10652 9024 10660 9033
rect 11057 9027 11115 9033
rect 11057 9024 11069 9027
rect 10652 8996 11069 9024
rect 10652 8987 10660 8996
rect 11057 8993 11069 8996
rect 11103 8993 11115 9027
rect 11057 8987 11115 8993
rect 10652 8984 10658 8987
rect 11146 8984 11152 9036
rect 11204 9024 11210 9036
rect 11330 9024 11336 9036
rect 11204 8996 11249 9024
rect 11291 8996 11336 9024
rect 11204 8984 11210 8996
rect 11330 8984 11336 8996
rect 11388 8984 11394 9036
rect 11790 9024 11796 9036
rect 11751 8996 11796 9024
rect 11790 8984 11796 8996
rect 11848 8984 11854 9036
rect 12268 9033 12296 9132
rect 12710 9120 12716 9132
rect 12768 9120 12774 9172
rect 12253 9027 12311 9033
rect 12253 8993 12265 9027
rect 12299 8993 12311 9027
rect 12894 9024 12900 9036
rect 12855 8996 12900 9024
rect 12253 8987 12311 8993
rect 12894 8984 12900 8996
rect 12952 9024 12958 9036
rect 13357 9027 13415 9033
rect 13357 9024 13369 9027
rect 12952 8996 13369 9024
rect 12952 8984 12958 8996
rect 13357 8993 13369 8996
rect 13403 8993 13415 9027
rect 13357 8987 13415 8993
rect 12345 8959 12403 8965
rect 12345 8956 12357 8959
rect 10300 8928 12357 8956
rect 9586 8919 9644 8925
rect 12345 8925 12357 8928
rect 12391 8925 12403 8959
rect 12345 8919 12403 8925
rect 7892 8860 8156 8888
rect 8481 8891 8539 8897
rect 7892 8848 7898 8860
rect 8481 8857 8493 8891
rect 8527 8888 8539 8891
rect 8754 8888 8760 8900
rect 8527 8860 8760 8888
rect 8527 8857 8539 8860
rect 8481 8851 8539 8857
rect 8754 8848 8760 8860
rect 8812 8848 8818 8900
rect 8938 8848 8944 8900
rect 8996 8888 9002 8900
rect 9600 8888 9628 8919
rect 11146 8888 11152 8900
rect 8996 8860 11152 8888
rect 8996 8848 9002 8860
rect 11146 8848 11152 8860
rect 11204 8848 11210 8900
rect 11974 8848 11980 8900
rect 12032 8888 12038 8900
rect 13173 8891 13231 8897
rect 13173 8888 13185 8891
rect 12032 8860 13185 8888
rect 12032 8848 12038 8860
rect 13173 8857 13185 8860
rect 13219 8857 13231 8891
rect 13173 8851 13231 8857
rect 6730 8820 6736 8832
rect 5644 8792 6736 8820
rect 4709 8783 4767 8789
rect 6730 8780 6736 8792
rect 6788 8820 6794 8832
rect 7098 8820 7104 8832
rect 6788 8792 7104 8820
rect 6788 8780 6794 8792
rect 7098 8780 7104 8792
rect 7156 8780 7162 8832
rect 8110 8780 8116 8832
rect 8168 8820 8174 8832
rect 9122 8820 9128 8832
rect 8168 8792 9128 8820
rect 8168 8780 8174 8792
rect 9122 8780 9128 8792
rect 9180 8820 9186 8832
rect 9490 8820 9496 8832
rect 9180 8792 9496 8820
rect 9180 8780 9186 8792
rect 9490 8780 9496 8792
rect 9548 8780 9554 8832
rect 9674 8780 9680 8832
rect 9732 8820 9738 8832
rect 9769 8823 9827 8829
rect 9769 8820 9781 8823
rect 9732 8792 9781 8820
rect 9732 8780 9738 8792
rect 9769 8789 9781 8792
rect 9815 8789 9827 8823
rect 9769 8783 9827 8789
rect 9858 8780 9864 8832
rect 9916 8820 9922 8832
rect 11241 8823 11299 8829
rect 11241 8820 11253 8823
rect 9916 8792 11253 8820
rect 9916 8780 9922 8792
rect 11241 8789 11253 8792
rect 11287 8789 11299 8823
rect 11241 8783 11299 8789
rect 1104 8730 13892 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 12246 8730
rect 12298 8678 12310 8730
rect 12362 8678 12374 8730
rect 12426 8678 12438 8730
rect 12490 8678 13892 8730
rect 1104 8656 13892 8678
rect 5350 8616 5356 8628
rect 5311 8588 5356 8616
rect 5350 8576 5356 8588
rect 5408 8576 5414 8628
rect 6086 8616 6092 8628
rect 6047 8588 6092 8616
rect 6086 8576 6092 8588
rect 6144 8576 6150 8628
rect 7098 8616 7104 8628
rect 7059 8588 7104 8616
rect 7098 8576 7104 8588
rect 7156 8576 7162 8628
rect 8662 8616 8668 8628
rect 8623 8588 8668 8616
rect 8662 8576 8668 8588
rect 8720 8576 8726 8628
rect 8754 8576 8760 8628
rect 8812 8616 8818 8628
rect 11330 8616 11336 8628
rect 8812 8588 11336 8616
rect 8812 8576 8818 8588
rect 11330 8576 11336 8588
rect 11388 8576 11394 8628
rect 3326 8508 3332 8560
rect 3384 8508 3390 8560
rect 5368 8548 5396 8576
rect 6917 8551 6975 8557
rect 6917 8548 6929 8551
rect 5368 8520 6929 8548
rect 6917 8517 6929 8520
rect 6963 8517 6975 8551
rect 6917 8511 6975 8517
rect 7926 8508 7932 8560
rect 7984 8548 7990 8560
rect 8202 8548 8208 8560
rect 7984 8520 8208 8548
rect 7984 8508 7990 8520
rect 8202 8508 8208 8520
rect 8260 8508 8266 8560
rect 9214 8508 9220 8560
rect 9272 8548 9278 8560
rect 10134 8548 10140 8560
rect 9272 8520 9536 8548
rect 9272 8508 9278 8520
rect 2038 8480 2044 8492
rect 1999 8452 2044 8480
rect 2038 8440 2044 8452
rect 2096 8440 2102 8492
rect 3344 8480 3372 8508
rect 6178 8480 6184 8492
rect 3344 8452 6184 8480
rect 1762 8412 1768 8424
rect 1723 8384 1768 8412
rect 1762 8372 1768 8384
rect 1820 8372 1826 8424
rect 2685 8415 2743 8421
rect 2685 8381 2697 8415
rect 2731 8412 2743 8415
rect 2866 8412 2872 8424
rect 2731 8384 2872 8412
rect 2731 8381 2743 8384
rect 2685 8375 2743 8381
rect 2866 8372 2872 8384
rect 2924 8372 2930 8424
rect 3344 8421 3372 8452
rect 6178 8440 6184 8452
rect 6236 8440 6242 8492
rect 7006 8480 7012 8492
rect 6919 8452 7012 8480
rect 7006 8440 7012 8452
rect 7064 8480 7070 8492
rect 9125 8483 9183 8489
rect 7064 8452 9076 8480
rect 7064 8440 7070 8452
rect 3329 8415 3387 8421
rect 3329 8381 3341 8415
rect 3375 8381 3387 8415
rect 3602 8412 3608 8424
rect 3563 8384 3608 8412
rect 3329 8375 3387 8381
rect 3602 8372 3608 8384
rect 3660 8372 3666 8424
rect 5810 8372 5816 8424
rect 5868 8412 5874 8424
rect 5905 8415 5963 8421
rect 5905 8412 5917 8415
rect 5868 8384 5917 8412
rect 5868 8372 5874 8384
rect 5905 8381 5917 8384
rect 5951 8381 5963 8415
rect 6822 8412 6828 8424
rect 6783 8384 6828 8412
rect 5905 8375 5963 8381
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 7193 8415 7251 8421
rect 7193 8381 7205 8415
rect 7239 8381 7251 8415
rect 7193 8375 7251 8381
rect 1854 8344 1860 8356
rect 1815 8316 1860 8344
rect 1854 8304 1860 8316
rect 1912 8304 1918 8356
rect 2406 8344 2412 8356
rect 2367 8316 2412 8344
rect 2406 8304 2412 8316
rect 2464 8304 2470 8356
rect 3881 8347 3939 8353
rect 3881 8313 3893 8347
rect 3927 8344 3939 8347
rect 4154 8344 4160 8356
rect 3927 8316 4160 8344
rect 3927 8313 3939 8316
rect 3881 8307 3939 8313
rect 4154 8304 4160 8316
rect 4212 8304 4218 8356
rect 5626 8344 5632 8356
rect 5106 8316 5632 8344
rect 5626 8304 5632 8316
rect 5684 8304 5690 8356
rect 7208 8344 7236 8375
rect 7558 8372 7564 8424
rect 7616 8412 7622 8424
rect 7653 8415 7711 8421
rect 7653 8412 7665 8415
rect 7616 8384 7665 8412
rect 7616 8372 7622 8384
rect 7653 8381 7665 8384
rect 7699 8381 7711 8415
rect 7653 8375 7711 8381
rect 7742 8372 7748 8424
rect 7800 8412 7806 8424
rect 8026 8415 8084 8421
rect 8026 8412 8038 8415
rect 7800 8384 8038 8412
rect 7800 8372 7806 8384
rect 8026 8381 8038 8384
rect 8072 8412 8084 8415
rect 8072 8384 8294 8412
rect 8072 8381 8084 8384
rect 8026 8375 8084 8381
rect 5736 8316 7236 8344
rect 1394 8276 1400 8288
rect 1355 8248 1400 8276
rect 1394 8236 1400 8248
rect 1452 8236 1458 8288
rect 4890 8236 4896 8288
rect 4948 8276 4954 8288
rect 5736 8276 5764 8316
rect 7282 8304 7288 8356
rect 7340 8344 7346 8356
rect 7837 8347 7895 8353
rect 7837 8344 7849 8347
rect 7340 8316 7849 8344
rect 7340 8304 7346 8316
rect 7837 8313 7849 8316
rect 7883 8313 7895 8347
rect 7837 8307 7895 8313
rect 7929 8347 7987 8353
rect 7929 8313 7941 8347
rect 7975 8344 7987 8347
rect 8110 8344 8116 8356
rect 7975 8316 8116 8344
rect 7975 8313 7987 8316
rect 7929 8307 7987 8313
rect 8110 8304 8116 8316
rect 8168 8304 8174 8356
rect 8266 8344 8294 8384
rect 8754 8372 8760 8424
rect 8812 8412 8818 8424
rect 8938 8412 8944 8424
rect 8812 8384 8857 8412
rect 8899 8384 8944 8412
rect 8812 8372 8818 8384
rect 8938 8372 8944 8384
rect 8996 8372 9002 8424
rect 9048 8412 9076 8452
rect 9125 8449 9137 8483
rect 9171 8480 9183 8483
rect 9306 8480 9312 8492
rect 9171 8452 9312 8480
rect 9171 8449 9183 8452
rect 9125 8443 9183 8449
rect 9306 8440 9312 8452
rect 9364 8440 9370 8492
rect 9508 8424 9536 8520
rect 9600 8520 10140 8548
rect 9217 8415 9275 8421
rect 9217 8412 9229 8415
rect 9048 8384 9229 8412
rect 9217 8381 9229 8384
rect 9263 8412 9275 8415
rect 9490 8412 9496 8424
rect 9263 8384 9352 8412
rect 9451 8384 9496 8412
rect 9263 8381 9275 8384
rect 9217 8375 9275 8381
rect 9125 8347 9183 8353
rect 9125 8344 9137 8347
rect 8266 8316 9137 8344
rect 9125 8313 9137 8316
rect 9171 8313 9183 8347
rect 9125 8307 9183 8313
rect 5902 8276 5908 8288
rect 4948 8248 5908 8276
rect 4948 8236 4954 8248
rect 5902 8236 5908 8248
rect 5960 8236 5966 8288
rect 6546 8276 6552 8288
rect 6507 8248 6552 8276
rect 6546 8236 6552 8248
rect 6604 8236 6610 8288
rect 9324 8276 9352 8384
rect 9490 8372 9496 8384
rect 9548 8372 9554 8424
rect 9600 8421 9628 8520
rect 10134 8508 10140 8520
rect 10192 8548 10198 8560
rect 10502 8548 10508 8560
rect 10192 8520 10272 8548
rect 10463 8520 10508 8548
rect 10192 8508 10198 8520
rect 9585 8415 9643 8421
rect 9585 8381 9597 8415
rect 9631 8381 9643 8415
rect 9585 8375 9643 8381
rect 9769 8415 9827 8421
rect 9769 8381 9781 8415
rect 9815 8412 9827 8415
rect 10042 8412 10048 8424
rect 9815 8384 10048 8412
rect 9815 8381 9827 8384
rect 9769 8375 9827 8381
rect 9398 8304 9404 8356
rect 9456 8344 9462 8356
rect 9600 8344 9628 8375
rect 10042 8372 10048 8384
rect 10100 8372 10106 8424
rect 10244 8412 10272 8520
rect 10502 8508 10508 8520
rect 10560 8508 10566 8560
rect 11790 8508 11796 8560
rect 11848 8548 11854 8560
rect 13081 8551 13139 8557
rect 13081 8548 13093 8551
rect 11848 8520 13093 8548
rect 11848 8508 11854 8520
rect 13081 8517 13093 8520
rect 13127 8517 13139 8551
rect 13081 8511 13139 8517
rect 10686 8440 10692 8492
rect 10744 8480 10750 8492
rect 12713 8483 12771 8489
rect 10744 8452 11008 8480
rect 10744 8440 10750 8452
rect 10321 8415 10379 8421
rect 10321 8412 10333 8415
rect 10244 8384 10333 8412
rect 10321 8381 10333 8384
rect 10367 8381 10379 8415
rect 10321 8375 10379 8381
rect 10505 8415 10563 8421
rect 10505 8381 10517 8415
rect 10551 8412 10563 8415
rect 10870 8412 10876 8424
rect 10551 8384 10876 8412
rect 10551 8381 10563 8384
rect 10505 8375 10563 8381
rect 10870 8372 10876 8384
rect 10928 8372 10934 8424
rect 10980 8421 11008 8452
rect 12713 8449 12725 8483
rect 12759 8480 12771 8483
rect 12802 8480 12808 8492
rect 12759 8452 12808 8480
rect 12759 8449 12771 8452
rect 12713 8443 12771 8449
rect 12802 8440 12808 8452
rect 12860 8440 12866 8492
rect 10965 8415 11023 8421
rect 10965 8381 10977 8415
rect 11011 8381 11023 8415
rect 10965 8375 11023 8381
rect 12437 8415 12495 8421
rect 12437 8381 12449 8415
rect 12483 8412 12495 8415
rect 12526 8412 12532 8424
rect 12483 8384 12532 8412
rect 12483 8381 12495 8384
rect 12437 8375 12495 8381
rect 12526 8372 12532 8384
rect 12584 8372 12590 8424
rect 12894 8372 12900 8424
rect 12952 8412 12958 8424
rect 13265 8415 13323 8421
rect 13265 8412 13277 8415
rect 12952 8384 13277 8412
rect 12952 8372 12958 8384
rect 13265 8381 13277 8384
rect 13311 8381 13323 8415
rect 13265 8375 13323 8381
rect 10134 8344 10140 8356
rect 9456 8316 9628 8344
rect 10095 8316 10140 8344
rect 9456 8304 9462 8316
rect 10134 8304 10140 8316
rect 10192 8304 10198 8356
rect 10226 8304 10232 8356
rect 10284 8344 10290 8356
rect 11057 8347 11115 8353
rect 11057 8344 11069 8347
rect 10284 8316 11069 8344
rect 10284 8304 10290 8316
rect 11057 8313 11069 8316
rect 11103 8313 11115 8347
rect 12618 8344 12624 8356
rect 11057 8307 11115 8313
rect 12544 8316 12624 8344
rect 9766 8276 9772 8288
rect 9324 8248 9772 8276
rect 9766 8236 9772 8248
rect 9824 8276 9830 8288
rect 10410 8276 10416 8288
rect 9824 8248 10416 8276
rect 9824 8236 9830 8248
rect 10410 8236 10416 8248
rect 10468 8236 10474 8288
rect 12066 8276 12072 8288
rect 12027 8248 12072 8276
rect 12066 8236 12072 8248
rect 12124 8236 12130 8288
rect 12544 8285 12572 8316
rect 12618 8304 12624 8316
rect 12676 8304 12682 8356
rect 12529 8279 12587 8285
rect 12529 8245 12541 8279
rect 12575 8245 12587 8279
rect 12529 8239 12587 8245
rect 1104 8186 13892 8208
rect 1104 8134 8246 8186
rect 8298 8134 8310 8186
rect 8362 8134 8374 8186
rect 8426 8134 8438 8186
rect 8490 8134 13892 8186
rect 1104 8112 13892 8134
rect 4154 8032 4160 8084
rect 4212 8072 4218 8084
rect 4709 8075 4767 8081
rect 4709 8072 4721 8075
rect 4212 8044 4721 8072
rect 4212 8032 4218 8044
rect 4709 8041 4721 8044
rect 4755 8041 4767 8075
rect 4709 8035 4767 8041
rect 4893 8075 4951 8081
rect 4893 8041 4905 8075
rect 4939 8072 4951 8075
rect 5445 8075 5503 8081
rect 5445 8072 5457 8075
rect 4939 8044 5457 8072
rect 4939 8041 4951 8044
rect 4893 8035 4951 8041
rect 5445 8041 5457 8044
rect 5491 8041 5503 8075
rect 5626 8072 5632 8084
rect 5587 8044 5632 8072
rect 5445 8035 5503 8041
rect 5626 8032 5632 8044
rect 5684 8032 5690 8084
rect 6178 8072 6184 8084
rect 6139 8044 6184 8072
rect 6178 8032 6184 8044
rect 6236 8032 6242 8084
rect 6549 8075 6607 8081
rect 6549 8041 6561 8075
rect 6595 8072 6607 8075
rect 6638 8072 6644 8084
rect 6595 8044 6644 8072
rect 6595 8041 6607 8044
rect 6549 8035 6607 8041
rect 6638 8032 6644 8044
rect 6696 8032 6702 8084
rect 9674 8072 9680 8084
rect 9416 8044 9680 8072
rect 3878 7964 3884 8016
rect 3936 8004 3942 8016
rect 4065 8007 4123 8013
rect 4065 8004 4077 8007
rect 3936 7976 4077 8004
rect 3936 7964 3942 7976
rect 4065 7973 4077 7976
rect 4111 7973 4123 8007
rect 4065 7967 4123 7973
rect 4818 7976 5580 8004
rect 1394 7896 1400 7948
rect 1452 7936 1458 7948
rect 1489 7939 1547 7945
rect 1489 7936 1501 7939
rect 1452 7908 1501 7936
rect 1452 7896 1458 7908
rect 1489 7905 1501 7908
rect 1535 7905 1547 7939
rect 1489 7899 1547 7905
rect 2406 7896 2412 7948
rect 2464 7936 2470 7948
rect 2961 7939 3019 7945
rect 2961 7936 2973 7939
rect 2464 7908 2973 7936
rect 2464 7896 2470 7908
rect 2961 7905 2973 7908
rect 3007 7905 3019 7939
rect 3326 7936 3332 7948
rect 3287 7908 3332 7936
rect 2961 7899 3019 7905
rect 2976 7868 3004 7899
rect 3326 7896 3332 7908
rect 3384 7936 3390 7948
rect 3970 7936 3976 7948
rect 3384 7908 3976 7936
rect 3384 7896 3390 7908
rect 3970 7896 3976 7908
rect 4028 7936 4034 7948
rect 4818 7936 4846 7976
rect 4028 7908 4846 7936
rect 4891 7939 4949 7945
rect 4028 7896 4034 7908
rect 4891 7905 4903 7939
rect 4937 7936 4949 7939
rect 5350 7936 5356 7948
rect 4937 7908 5356 7936
rect 4937 7905 4949 7908
rect 4891 7899 4949 7905
rect 5350 7896 5356 7908
rect 5408 7936 5414 7948
rect 5552 7936 5580 7976
rect 7742 7964 7748 8016
rect 7800 8004 7806 8016
rect 9416 8013 9444 8044
rect 9674 8032 9680 8044
rect 9732 8032 9738 8084
rect 9769 8075 9827 8081
rect 9769 8041 9781 8075
rect 9815 8072 9827 8075
rect 10134 8072 10140 8084
rect 9815 8044 10140 8072
rect 9815 8041 9827 8044
rect 9769 8035 9827 8041
rect 10134 8032 10140 8044
rect 10192 8032 10198 8084
rect 10410 8032 10416 8084
rect 10468 8072 10474 8084
rect 11977 8075 12035 8081
rect 11977 8072 11989 8075
rect 10468 8044 11989 8072
rect 10468 8032 10474 8044
rect 11977 8041 11989 8044
rect 12023 8041 12035 8075
rect 11977 8035 12035 8041
rect 7929 8007 7987 8013
rect 7929 8004 7941 8007
rect 7800 7976 7941 8004
rect 7800 7964 7806 7976
rect 7929 7973 7941 7976
rect 7975 7973 7987 8007
rect 7929 7967 7987 7973
rect 9401 8007 9459 8013
rect 9401 7973 9413 8007
rect 9447 7973 9459 8007
rect 9401 7967 9459 7973
rect 9493 8007 9551 8013
rect 9493 7973 9505 8007
rect 9539 8004 9551 8007
rect 10226 8004 10232 8016
rect 9539 7976 10232 8004
rect 9539 7973 9551 7976
rect 9493 7967 9551 7973
rect 10226 7964 10232 7976
rect 10284 7964 10290 8016
rect 10502 8004 10508 8016
rect 10463 7976 10508 8004
rect 10502 7964 10508 7976
rect 10560 7964 10566 8016
rect 11790 8004 11796 8016
rect 11730 7976 11796 8004
rect 11790 7964 11796 7976
rect 11848 7964 11854 8016
rect 13081 8007 13139 8013
rect 13081 7973 13093 8007
rect 13127 8004 13139 8007
rect 13354 8004 13360 8016
rect 13127 7976 13360 8004
rect 13127 7973 13139 7976
rect 13081 7967 13139 7973
rect 13354 7964 13360 7976
rect 13412 7964 13418 8016
rect 5810 7936 5816 7948
rect 5408 7908 5453 7936
rect 5552 7908 5816 7936
rect 5408 7896 5414 7908
rect 5810 7896 5816 7908
rect 5868 7896 5874 7948
rect 6641 7939 6699 7945
rect 6641 7905 6653 7939
rect 6687 7936 6699 7939
rect 6914 7936 6920 7948
rect 6687 7908 6920 7936
rect 6687 7905 6699 7908
rect 6641 7899 6699 7905
rect 6914 7896 6920 7908
rect 6972 7896 6978 7948
rect 7190 7936 7196 7948
rect 7151 7908 7196 7936
rect 7190 7896 7196 7908
rect 7248 7936 7254 7948
rect 7374 7936 7380 7948
rect 7248 7908 7380 7936
rect 7248 7896 7254 7908
rect 7374 7896 7380 7908
rect 7432 7936 7438 7948
rect 8021 7939 8079 7945
rect 8021 7936 8033 7939
rect 7432 7908 8033 7936
rect 7432 7896 7438 7908
rect 8021 7905 8033 7908
rect 8067 7936 8079 7939
rect 8110 7936 8116 7948
rect 8067 7908 8116 7936
rect 8067 7905 8079 7908
rect 8021 7899 8079 7905
rect 8110 7896 8116 7908
rect 8168 7896 8174 7948
rect 9122 7936 9128 7948
rect 9083 7908 9128 7936
rect 9122 7896 9128 7908
rect 9180 7896 9186 7948
rect 9273 7939 9331 7945
rect 9273 7905 9285 7939
rect 9319 7936 9331 7939
rect 9631 7939 9689 7945
rect 9319 7905 9352 7936
rect 9273 7899 9352 7905
rect 9631 7905 9643 7939
rect 9677 7936 9689 7939
rect 10042 7936 10048 7948
rect 9677 7908 10048 7936
rect 9677 7905 9689 7908
rect 9631 7899 9689 7905
rect 3881 7871 3939 7877
rect 3881 7868 3893 7871
rect 2976 7840 3893 7868
rect 3881 7837 3893 7840
rect 3927 7837 3939 7871
rect 6822 7868 6828 7880
rect 6783 7840 6828 7868
rect 3881 7831 3939 7837
rect 6822 7828 6828 7840
rect 6880 7828 6886 7880
rect 7834 7868 7840 7880
rect 7795 7840 7840 7868
rect 7834 7828 7840 7840
rect 7892 7828 7898 7880
rect 2958 7800 2964 7812
rect 2919 7772 2964 7800
rect 2958 7760 2964 7772
rect 3016 7760 3022 7812
rect 3513 7803 3571 7809
rect 3513 7769 3525 7803
rect 3559 7800 3571 7803
rect 6362 7800 6368 7812
rect 3559 7772 6368 7800
rect 3559 7769 3571 7772
rect 3513 7763 3571 7769
rect 6362 7760 6368 7772
rect 6420 7760 6426 7812
rect 5261 7735 5319 7741
rect 5261 7701 5273 7735
rect 5307 7732 5319 7735
rect 5445 7735 5503 7741
rect 5445 7732 5457 7735
rect 5307 7704 5457 7732
rect 5307 7701 5319 7704
rect 5261 7695 5319 7701
rect 5445 7701 5457 7704
rect 5491 7732 5503 7735
rect 5902 7732 5908 7744
rect 5491 7704 5908 7732
rect 5491 7701 5503 7704
rect 5445 7695 5503 7701
rect 5902 7692 5908 7704
rect 5960 7692 5966 7744
rect 7282 7732 7288 7744
rect 7243 7704 7288 7732
rect 7282 7692 7288 7704
rect 7340 7692 7346 7744
rect 8018 7692 8024 7744
rect 8076 7732 8082 7744
rect 8389 7735 8447 7741
rect 8389 7732 8401 7735
rect 8076 7704 8401 7732
rect 8076 7692 8082 7704
rect 8389 7701 8401 7704
rect 8435 7701 8447 7735
rect 9324 7732 9352 7899
rect 10042 7896 10048 7908
rect 10100 7896 10106 7948
rect 12066 7896 12072 7948
rect 12124 7936 12130 7948
rect 12345 7939 12403 7945
rect 12345 7936 12357 7939
rect 12124 7908 12357 7936
rect 12124 7896 12130 7908
rect 12345 7905 12357 7908
rect 12391 7905 12403 7939
rect 13262 7936 13268 7948
rect 13223 7908 13268 7936
rect 12345 7899 12403 7905
rect 13262 7896 13268 7908
rect 13320 7896 13326 7948
rect 10226 7868 10232 7880
rect 10187 7840 10232 7868
rect 10226 7828 10232 7840
rect 10284 7868 10290 7880
rect 10594 7868 10600 7880
rect 10284 7840 10600 7868
rect 10284 7828 10290 7840
rect 10594 7828 10600 7840
rect 10652 7828 10658 7880
rect 10870 7732 10876 7744
rect 9324 7704 10876 7732
rect 8389 7695 8447 7701
rect 10870 7692 10876 7704
rect 10928 7692 10934 7744
rect 1104 7642 13892 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 12246 7642
rect 12298 7590 12310 7642
rect 12362 7590 12374 7642
rect 12426 7590 12438 7642
rect 12490 7590 13892 7642
rect 1104 7568 13892 7590
rect 5810 7528 5816 7540
rect 5368 7500 5816 7528
rect 5368 7469 5396 7500
rect 5810 7488 5816 7500
rect 5868 7528 5874 7540
rect 7650 7528 7656 7540
rect 5868 7500 7656 7528
rect 5868 7488 5874 7500
rect 7650 7488 7656 7500
rect 7708 7488 7714 7540
rect 9122 7528 9128 7540
rect 7760 7500 9128 7528
rect 5353 7463 5411 7469
rect 5353 7429 5365 7463
rect 5399 7429 5411 7463
rect 5353 7423 5411 7429
rect 6822 7420 6828 7472
rect 6880 7420 6886 7472
rect 1394 7352 1400 7404
rect 1452 7392 1458 7404
rect 1949 7395 2007 7401
rect 1949 7392 1961 7395
rect 1452 7364 1961 7392
rect 1452 7352 1458 7364
rect 1949 7361 1961 7364
rect 1995 7361 2007 7395
rect 1949 7355 2007 7361
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7392 2559 7395
rect 2774 7392 2780 7404
rect 2547 7364 2780 7392
rect 2547 7361 2559 7364
rect 2501 7355 2559 7361
rect 2774 7352 2780 7364
rect 2832 7352 2838 7404
rect 5258 7392 5264 7404
rect 5219 7364 5264 7392
rect 5258 7352 5264 7364
rect 5316 7352 5322 7404
rect 5442 7352 5448 7404
rect 5500 7392 5506 7404
rect 6840 7392 6868 7420
rect 7009 7395 7067 7401
rect 7009 7392 7021 7395
rect 5500 7364 7021 7392
rect 5500 7352 5506 7364
rect 7009 7361 7021 7364
rect 7055 7361 7067 7395
rect 7009 7355 7067 7361
rect 1489 7327 1547 7333
rect 1489 7293 1501 7327
rect 1535 7293 1547 7327
rect 1489 7287 1547 7293
rect 2409 7327 2467 7333
rect 2409 7293 2421 7327
rect 2455 7324 2467 7327
rect 2958 7324 2964 7336
rect 2455 7296 2964 7324
rect 2455 7293 2467 7296
rect 2409 7287 2467 7293
rect 1504 7256 1532 7287
rect 2958 7284 2964 7296
rect 3016 7284 3022 7336
rect 3326 7284 3332 7336
rect 3384 7324 3390 7336
rect 3421 7327 3479 7333
rect 3421 7324 3433 7327
rect 3384 7296 3433 7324
rect 3384 7284 3390 7296
rect 3421 7293 3433 7296
rect 3467 7293 3479 7327
rect 3421 7287 3479 7293
rect 2498 7256 2504 7268
rect 1504 7228 2504 7256
rect 2498 7216 2504 7228
rect 2556 7256 2562 7268
rect 2777 7259 2835 7265
rect 2777 7256 2789 7259
rect 2556 7228 2789 7256
rect 2556 7216 2562 7228
rect 2777 7225 2789 7228
rect 2823 7225 2835 7259
rect 3436 7256 3464 7287
rect 3510 7284 3516 7336
rect 3568 7324 3574 7336
rect 3881 7327 3939 7333
rect 3881 7324 3893 7327
rect 3568 7296 3893 7324
rect 3568 7284 3574 7296
rect 3881 7293 3893 7296
rect 3927 7293 3939 7327
rect 3881 7287 3939 7293
rect 4338 7284 4344 7336
rect 4396 7324 4402 7336
rect 5813 7327 5871 7333
rect 5813 7324 5825 7327
rect 4396 7296 5825 7324
rect 4396 7284 4402 7296
rect 5813 7293 5825 7296
rect 5859 7293 5871 7327
rect 5813 7287 5871 7293
rect 3786 7256 3792 7268
rect 3436 7228 3792 7256
rect 2777 7219 2835 7225
rect 3786 7216 3792 7228
rect 3844 7216 3850 7268
rect 4522 7256 4528 7268
rect 4483 7228 4528 7256
rect 4522 7216 4528 7228
rect 4580 7216 4586 7268
rect 4801 7259 4859 7265
rect 4801 7225 4813 7259
rect 4847 7256 4859 7259
rect 5074 7256 5080 7268
rect 4847 7228 5080 7256
rect 4847 7225 4859 7228
rect 4801 7219 4859 7225
rect 5074 7216 5080 7228
rect 5132 7256 5138 7268
rect 5626 7256 5632 7268
rect 5132 7228 5632 7256
rect 5132 7216 5138 7228
rect 5626 7216 5632 7228
rect 5684 7216 5690 7268
rect 1670 7188 1676 7200
rect 1631 7160 1676 7188
rect 1670 7148 1676 7160
rect 1728 7148 1734 7200
rect 3605 7191 3663 7197
rect 3605 7157 3617 7191
rect 3651 7188 3663 7191
rect 4614 7188 4620 7200
rect 3651 7160 4620 7188
rect 3651 7157 3663 7160
rect 3605 7151 3663 7157
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 5828 7188 5856 7287
rect 6546 7284 6552 7336
rect 6604 7324 6610 7336
rect 7760 7333 7788 7500
rect 9122 7488 9128 7500
rect 9180 7488 9186 7540
rect 10137 7531 10195 7537
rect 10137 7528 10149 7531
rect 9232 7500 10149 7528
rect 8110 7460 8116 7472
rect 8036 7432 8116 7460
rect 8036 7401 8064 7432
rect 8110 7420 8116 7432
rect 8168 7420 8174 7472
rect 8202 7420 8208 7472
rect 8260 7460 8266 7472
rect 8260 7432 8340 7460
rect 8260 7420 8266 7432
rect 8312 7401 8340 7432
rect 8004 7395 8064 7401
rect 8004 7361 8016 7395
rect 8050 7364 8064 7395
rect 8297 7395 8355 7401
rect 8050 7361 8062 7364
rect 8004 7355 8062 7361
rect 8297 7361 8309 7395
rect 8343 7361 8355 7395
rect 8297 7355 8355 7361
rect 6825 7327 6883 7333
rect 6825 7324 6837 7327
rect 6604 7296 6837 7324
rect 6604 7284 6610 7296
rect 6825 7293 6837 7296
rect 6871 7293 6883 7327
rect 7745 7327 7803 7333
rect 7745 7324 7757 7327
rect 6825 7287 6883 7293
rect 7300 7296 7757 7324
rect 6730 7216 6736 7268
rect 6788 7256 6794 7268
rect 7300 7256 7328 7296
rect 7745 7293 7757 7296
rect 7791 7293 7803 7327
rect 8082 7327 8140 7333
rect 8082 7324 8094 7327
rect 7745 7287 7803 7293
rect 7852 7296 8094 7324
rect 6788 7228 7328 7256
rect 6788 7216 6794 7228
rect 7374 7216 7380 7268
rect 7432 7256 7438 7268
rect 7561 7259 7619 7265
rect 7561 7256 7573 7259
rect 7432 7228 7573 7256
rect 7432 7216 7438 7228
rect 7561 7225 7573 7228
rect 7607 7225 7619 7259
rect 7561 7219 7619 7225
rect 7650 7216 7656 7268
rect 7708 7256 7714 7268
rect 7852 7256 7880 7296
rect 8082 7293 8094 7296
rect 8128 7293 8140 7327
rect 8082 7287 8140 7293
rect 9030 7284 9036 7336
rect 9088 7324 9094 7336
rect 9232 7333 9260 7500
rect 10137 7497 10149 7500
rect 10183 7497 10195 7531
rect 10137 7491 10195 7497
rect 10870 7488 10876 7540
rect 10928 7528 10934 7540
rect 12989 7531 13047 7537
rect 12989 7528 13001 7531
rect 10928 7500 13001 7528
rect 10928 7488 10934 7500
rect 12989 7497 13001 7500
rect 13035 7497 13047 7531
rect 12989 7491 13047 7497
rect 9490 7460 9496 7472
rect 9451 7432 9496 7460
rect 9490 7420 9496 7432
rect 9548 7420 9554 7472
rect 12529 7463 12587 7469
rect 12529 7429 12541 7463
rect 12575 7460 12587 7463
rect 13354 7460 13360 7472
rect 12575 7432 13360 7460
rect 12575 7429 12587 7432
rect 12529 7423 12587 7429
rect 13354 7420 13360 7432
rect 13412 7420 13418 7472
rect 9950 7352 9956 7404
rect 10008 7392 10014 7404
rect 10778 7392 10784 7404
rect 10008 7364 10364 7392
rect 10739 7364 10784 7392
rect 10008 7352 10014 7364
rect 9217 7327 9275 7333
rect 9217 7324 9229 7327
rect 9088 7296 9229 7324
rect 9088 7284 9094 7296
rect 9217 7293 9229 7296
rect 9263 7293 9275 7327
rect 9217 7287 9275 7293
rect 9309 7327 9367 7333
rect 9309 7293 9321 7327
rect 9355 7293 9367 7327
rect 9309 7287 9367 7293
rect 9585 7327 9643 7333
rect 9585 7293 9597 7327
rect 9631 7324 9643 7327
rect 9766 7324 9772 7336
rect 9631 7296 9772 7324
rect 9631 7293 9643 7296
rect 9585 7287 9643 7293
rect 9324 7256 9352 7287
rect 9766 7284 9772 7296
rect 9824 7324 9830 7336
rect 10336 7333 10364 7364
rect 10778 7352 10784 7364
rect 10836 7352 10842 7404
rect 11333 7395 11391 7401
rect 11333 7361 11345 7395
rect 11379 7392 11391 7395
rect 12621 7395 12679 7401
rect 11379 7364 12434 7392
rect 11379 7361 11391 7364
rect 11333 7355 11391 7361
rect 12406 7336 12434 7364
rect 12621 7361 12633 7395
rect 12667 7392 12679 7395
rect 12986 7392 12992 7404
rect 12667 7364 12992 7392
rect 12667 7361 12679 7364
rect 12621 7355 12679 7361
rect 12986 7352 12992 7364
rect 13044 7352 13050 7404
rect 10137 7327 10195 7333
rect 10137 7324 10149 7327
rect 9824 7296 10149 7324
rect 9824 7284 9830 7296
rect 10137 7293 10149 7296
rect 10183 7293 10195 7327
rect 10137 7287 10195 7293
rect 10321 7327 10379 7333
rect 10321 7293 10333 7327
rect 10367 7293 10379 7327
rect 12066 7324 12072 7336
rect 12027 7296 12072 7324
rect 10321 7287 10379 7293
rect 12066 7284 12072 7296
rect 12124 7284 12130 7336
rect 12406 7296 12440 7336
rect 12434 7284 12440 7296
rect 12492 7284 12498 7336
rect 12897 7327 12955 7333
rect 12897 7293 12909 7327
rect 12943 7293 12955 7327
rect 12897 7287 12955 7293
rect 9858 7256 9864 7268
rect 7708 7228 7880 7256
rect 7944 7228 9260 7256
rect 9324 7228 9864 7256
rect 7708 7216 7714 7228
rect 6457 7191 6515 7197
rect 6457 7188 6469 7191
rect 5828 7160 6469 7188
rect 6457 7157 6469 7160
rect 6503 7157 6515 7191
rect 6457 7151 6515 7157
rect 6917 7191 6975 7197
rect 6917 7157 6929 7191
rect 6963 7188 6975 7191
rect 7944 7188 7972 7228
rect 6963 7160 7972 7188
rect 8205 7191 8263 7197
rect 6963 7157 6975 7160
rect 6917 7151 6975 7157
rect 8205 7157 8217 7191
rect 8251 7188 8263 7191
rect 8662 7188 8668 7200
rect 8251 7160 8668 7188
rect 8251 7157 8263 7160
rect 8205 7151 8263 7157
rect 8662 7148 8668 7160
rect 8720 7148 8726 7200
rect 8754 7148 8760 7200
rect 8812 7188 8818 7200
rect 9033 7191 9091 7197
rect 9033 7188 9045 7191
rect 8812 7160 9045 7188
rect 8812 7148 8818 7160
rect 9033 7157 9045 7160
rect 9079 7157 9091 7191
rect 9232 7188 9260 7228
rect 9858 7216 9864 7228
rect 9916 7216 9922 7268
rect 11238 7256 11244 7268
rect 11199 7228 11244 7256
rect 11238 7216 11244 7228
rect 11296 7216 11302 7268
rect 9674 7188 9680 7200
rect 9232 7160 9680 7188
rect 9033 7151 9091 7157
rect 9674 7148 9680 7160
rect 9732 7148 9738 7200
rect 9950 7188 9956 7200
rect 9911 7160 9956 7188
rect 9950 7148 9956 7160
rect 10008 7148 10014 7200
rect 10042 7148 10048 7200
rect 10100 7188 10106 7200
rect 12912 7188 12940 7287
rect 10100 7160 12940 7188
rect 10100 7148 10106 7160
rect 1104 7098 13892 7120
rect 1104 7046 8246 7098
rect 8298 7046 8310 7098
rect 8362 7046 8374 7098
rect 8426 7046 8438 7098
rect 8490 7046 13892 7098
rect 1104 7024 13892 7046
rect 3145 6987 3203 6993
rect 3145 6953 3157 6987
rect 3191 6984 3203 6987
rect 4062 6984 4068 6996
rect 3191 6956 4068 6984
rect 3191 6953 3203 6956
rect 3145 6947 3203 6953
rect 4062 6944 4068 6956
rect 4120 6944 4126 6996
rect 7006 6944 7012 6996
rect 7064 6984 7070 6996
rect 7834 6984 7840 6996
rect 7064 6956 7840 6984
rect 7064 6944 7070 6956
rect 7834 6944 7840 6956
rect 7892 6984 7898 6996
rect 8754 6984 8760 6996
rect 7892 6956 8760 6984
rect 7892 6944 7898 6956
rect 2498 6916 2504 6928
rect 2459 6888 2504 6916
rect 2498 6876 2504 6888
rect 2556 6876 2562 6928
rect 7466 6876 7472 6928
rect 7524 6916 7530 6928
rect 8496 6925 8524 6956
rect 8754 6944 8760 6956
rect 8812 6944 8818 6996
rect 8481 6919 8539 6925
rect 7524 6888 8064 6916
rect 7524 6876 7530 6888
rect 1394 6808 1400 6860
rect 1452 6848 1458 6860
rect 1581 6851 1639 6857
rect 1581 6848 1593 6851
rect 1452 6820 1593 6848
rect 1452 6808 1458 6820
rect 1581 6817 1593 6820
rect 1627 6817 1639 6851
rect 1581 6811 1639 6817
rect 2130 6808 2136 6860
rect 2188 6848 2194 6860
rect 2225 6851 2283 6857
rect 2225 6848 2237 6851
rect 2188 6820 2237 6848
rect 2188 6808 2194 6820
rect 2225 6817 2237 6820
rect 2271 6817 2283 6851
rect 2225 6811 2283 6817
rect 2774 6808 2780 6860
rect 2832 6848 2838 6860
rect 3053 6851 3111 6857
rect 3053 6848 3065 6851
rect 2832 6820 3065 6848
rect 2832 6808 2838 6820
rect 3053 6817 3065 6820
rect 3099 6817 3111 6851
rect 3878 6848 3884 6860
rect 3839 6820 3884 6848
rect 3053 6811 3111 6817
rect 3878 6808 3884 6820
rect 3936 6808 3942 6860
rect 4338 6848 4344 6860
rect 4299 6820 4344 6848
rect 4338 6808 4344 6820
rect 4396 6808 4402 6860
rect 5626 6808 5632 6860
rect 5684 6848 5690 6860
rect 5813 6851 5871 6857
rect 5813 6848 5825 6851
rect 5684 6820 5825 6848
rect 5684 6808 5690 6820
rect 5813 6817 5825 6820
rect 5859 6848 5871 6851
rect 5997 6851 6055 6857
rect 5997 6848 6009 6851
rect 5859 6820 6009 6848
rect 5859 6817 5871 6820
rect 5813 6811 5871 6817
rect 5997 6817 6009 6820
rect 6043 6817 6055 6851
rect 5997 6811 6055 6817
rect 6178 6808 6184 6860
rect 6236 6848 6242 6860
rect 6454 6848 6460 6860
rect 6236 6820 6460 6848
rect 6236 6808 6242 6820
rect 6454 6808 6460 6820
rect 6512 6808 6518 6860
rect 8036 6857 8064 6888
rect 8481 6885 8493 6919
rect 8527 6885 8539 6919
rect 11238 6916 11244 6928
rect 8481 6879 8539 6885
rect 8588 6888 9260 6916
rect 11199 6888 11244 6916
rect 8021 6851 8079 6857
rect 2038 6740 2044 6792
rect 2096 6780 2102 6792
rect 2640 6784 2698 6790
rect 2640 6780 2652 6784
rect 2096 6752 2652 6780
rect 2096 6740 2102 6752
rect 2640 6750 2652 6752
rect 2686 6780 2698 6784
rect 2961 6783 3019 6789
rect 2961 6780 2973 6783
rect 2686 6752 2973 6780
rect 2686 6750 2698 6752
rect 2640 6744 2698 6750
rect 2961 6749 2973 6752
rect 3007 6780 3019 6783
rect 6656 6780 6684 6834
rect 8021 6817 8033 6851
rect 8067 6817 8079 6851
rect 8021 6811 8079 6817
rect 8202 6808 8208 6860
rect 8260 6848 8266 6860
rect 8297 6851 8355 6857
rect 8297 6848 8309 6851
rect 8260 6820 8309 6848
rect 8260 6808 8266 6820
rect 8297 6817 8309 6820
rect 8343 6817 8355 6851
rect 8297 6811 8355 6817
rect 8588 6780 8616 6888
rect 8754 6808 8760 6860
rect 8812 6848 8818 6860
rect 9125 6851 9183 6857
rect 9125 6848 9137 6851
rect 8812 6820 9137 6848
rect 8812 6808 8818 6820
rect 9125 6817 9137 6820
rect 9171 6817 9183 6851
rect 9232 6848 9260 6888
rect 11238 6876 11244 6888
rect 11296 6876 11302 6928
rect 12066 6876 12072 6928
rect 12124 6876 12130 6928
rect 9677 6851 9735 6857
rect 9232 6820 9536 6848
rect 9125 6811 9183 6817
rect 3007 6752 4016 6780
rect 3007 6749 3019 6752
rect 2961 6743 3019 6749
rect 3510 6644 3516 6656
rect 3471 6616 3516 6644
rect 3510 6604 3516 6616
rect 3568 6604 3574 6656
rect 3988 6644 4016 6752
rect 4080 6752 6684 6780
rect 6748 6752 8616 6780
rect 4080 6721 4108 6752
rect 4065 6715 4123 6721
rect 4065 6681 4077 6715
rect 4111 6681 4123 6715
rect 5810 6712 5816 6724
rect 5771 6684 5816 6712
rect 4065 6675 4123 6681
rect 5810 6672 5816 6684
rect 5868 6672 5874 6724
rect 5997 6715 6055 6721
rect 5997 6681 6009 6715
rect 6043 6712 6055 6715
rect 6748 6712 6776 6752
rect 8662 6740 8668 6792
rect 8720 6780 8726 6792
rect 9398 6780 9404 6792
rect 8720 6752 9404 6780
rect 8720 6740 8726 6752
rect 9398 6740 9404 6752
rect 9456 6740 9462 6792
rect 9508 6780 9536 6820
rect 9677 6817 9689 6851
rect 9723 6848 9735 6851
rect 10778 6848 10784 6860
rect 9723 6820 10784 6848
rect 9723 6817 9735 6820
rect 9677 6811 9735 6817
rect 10778 6808 10784 6820
rect 10836 6808 10842 6860
rect 11149 6851 11207 6857
rect 11149 6817 11161 6851
rect 11195 6817 11207 6851
rect 11149 6811 11207 6817
rect 10962 6780 10968 6792
rect 9508 6752 10968 6780
rect 10962 6740 10968 6752
rect 11020 6740 11026 6792
rect 11164 6780 11192 6811
rect 12710 6780 12716 6792
rect 11164 6752 12716 6780
rect 12710 6740 12716 6752
rect 12768 6740 12774 6792
rect 13078 6780 13084 6792
rect 13039 6752 13084 6780
rect 13078 6740 13084 6752
rect 13136 6740 13142 6792
rect 13357 6783 13415 6789
rect 13357 6749 13369 6783
rect 13403 6749 13415 6783
rect 13357 6743 13415 6749
rect 6043 6684 6776 6712
rect 6043 6681 6055 6684
rect 5997 6675 6055 6681
rect 8478 6672 8484 6724
rect 8536 6712 8542 6724
rect 8536 6684 8616 6712
rect 8536 6672 8542 6684
rect 5442 6644 5448 6656
rect 3988 6616 5448 6644
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 6273 6647 6331 6653
rect 6273 6613 6285 6647
rect 6319 6644 6331 6647
rect 7190 6644 7196 6656
rect 6319 6616 7196 6644
rect 6319 6613 6331 6616
rect 6273 6607 6331 6613
rect 7190 6604 7196 6616
rect 7248 6604 7254 6656
rect 7374 6604 7380 6656
rect 7432 6644 7438 6656
rect 8588 6653 8616 6684
rect 9122 6672 9128 6724
rect 9180 6712 9186 6724
rect 11422 6712 11428 6724
rect 9180 6684 11428 6712
rect 9180 6672 9186 6684
rect 11422 6672 11428 6684
rect 11480 6672 11486 6724
rect 11514 6672 11520 6724
rect 11572 6712 11578 6724
rect 11572 6684 11836 6712
rect 11572 6672 11578 6684
rect 7757 6647 7815 6653
rect 7757 6644 7769 6647
rect 7432 6616 7769 6644
rect 7432 6604 7438 6616
rect 7757 6613 7769 6616
rect 7803 6613 7815 6647
rect 7757 6607 7815 6613
rect 8573 6647 8631 6653
rect 8573 6613 8585 6647
rect 8619 6613 8631 6647
rect 8573 6607 8631 6613
rect 9030 6604 9036 6656
rect 9088 6644 9094 6656
rect 9217 6647 9275 6653
rect 9217 6644 9229 6647
rect 9088 6616 9229 6644
rect 9088 6604 9094 6616
rect 9217 6613 9229 6616
rect 9263 6613 9275 6647
rect 9217 6607 9275 6613
rect 9490 6604 9496 6656
rect 9548 6644 9554 6656
rect 10042 6644 10048 6656
rect 9548 6616 10048 6644
rect 9548 6604 9554 6616
rect 10042 6604 10048 6616
rect 10100 6644 10106 6656
rect 10502 6644 10508 6656
rect 10100 6616 10508 6644
rect 10100 6604 10106 6616
rect 10502 6604 10508 6616
rect 10560 6604 10566 6656
rect 11609 6647 11667 6653
rect 11609 6613 11621 6647
rect 11655 6644 11667 6647
rect 11698 6644 11704 6656
rect 11655 6616 11704 6644
rect 11655 6613 11667 6616
rect 11609 6607 11667 6613
rect 11698 6604 11704 6616
rect 11756 6604 11762 6656
rect 11808 6644 11836 6684
rect 13372 6644 13400 6743
rect 11808 6616 13400 6644
rect 1104 6554 13892 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 12246 6554
rect 12298 6502 12310 6554
rect 12362 6502 12374 6554
rect 12426 6502 12438 6554
rect 12490 6502 13892 6554
rect 1104 6480 13892 6502
rect 7009 6443 7067 6449
rect 7009 6409 7021 6443
rect 7055 6440 7067 6443
rect 8110 6440 8116 6452
rect 7055 6412 8116 6440
rect 7055 6409 7067 6412
rect 7009 6403 7067 6409
rect 8110 6400 8116 6412
rect 8168 6400 8174 6452
rect 10321 6443 10379 6449
rect 10321 6440 10333 6443
rect 8956 6412 10333 6440
rect 1857 6375 1915 6381
rect 1857 6341 1869 6375
rect 1903 6372 1915 6375
rect 2130 6372 2136 6384
rect 1903 6344 2136 6372
rect 1903 6341 1915 6344
rect 1857 6335 1915 6341
rect 2130 6332 2136 6344
rect 2188 6332 2194 6384
rect 2501 6375 2559 6381
rect 2501 6341 2513 6375
rect 2547 6372 2559 6375
rect 2866 6372 2872 6384
rect 2547 6344 2872 6372
rect 2547 6341 2559 6344
rect 2501 6335 2559 6341
rect 2866 6332 2872 6344
rect 2924 6332 2930 6384
rect 4525 6375 4583 6381
rect 4525 6341 4537 6375
rect 4571 6372 4583 6375
rect 5810 6372 5816 6384
rect 4571 6344 5816 6372
rect 4571 6341 4583 6344
rect 4525 6335 4583 6341
rect 5810 6332 5816 6344
rect 5868 6332 5874 6384
rect 5902 6332 5908 6384
rect 5960 6372 5966 6384
rect 7377 6375 7435 6381
rect 7377 6372 7389 6375
rect 5960 6344 7389 6372
rect 5960 6332 5966 6344
rect 7377 6341 7389 6344
rect 7423 6341 7435 6375
rect 7377 6335 7435 6341
rect 7558 6332 7564 6384
rect 7616 6332 7622 6384
rect 7650 6332 7656 6384
rect 7708 6372 7714 6384
rect 7708 6344 7880 6372
rect 7708 6332 7714 6344
rect 1394 6304 1400 6316
rect 1355 6276 1400 6304
rect 1394 6264 1400 6276
rect 1452 6264 1458 6316
rect 1670 6264 1676 6316
rect 1728 6304 1734 6316
rect 1949 6307 2007 6313
rect 1949 6304 1961 6307
rect 1728 6276 1961 6304
rect 1728 6264 1734 6276
rect 1949 6273 1961 6276
rect 1995 6273 2007 6307
rect 3878 6304 3884 6316
rect 1949 6267 2007 6273
rect 2332 6276 3884 6304
rect 1578 6196 1584 6248
rect 1636 6236 1642 6248
rect 2332 6236 2360 6276
rect 3878 6264 3884 6276
rect 3936 6304 3942 6316
rect 5258 6304 5264 6316
rect 3936 6276 4384 6304
rect 5219 6276 5264 6304
rect 3936 6264 3942 6276
rect 2498 6236 2504 6248
rect 1636 6208 2360 6236
rect 2459 6208 2504 6236
rect 1636 6196 1642 6208
rect 2498 6196 2504 6208
rect 2556 6196 2562 6248
rect 4356 6245 4384 6276
rect 5258 6264 5264 6276
rect 5316 6264 5322 6316
rect 5442 6304 5448 6316
rect 5403 6276 5448 6304
rect 5442 6264 5448 6276
rect 5500 6264 5506 6316
rect 7576 6304 7604 6332
rect 7852 6304 7880 6344
rect 7926 6332 7932 6384
rect 7984 6372 7990 6384
rect 8202 6372 8208 6384
rect 7984 6344 8208 6372
rect 7984 6332 7990 6344
rect 8202 6332 8208 6344
rect 8260 6332 8266 6384
rect 6104 6276 7788 6304
rect 3789 6239 3847 6245
rect 3789 6205 3801 6239
rect 3835 6205 3847 6239
rect 3789 6199 3847 6205
rect 4341 6239 4399 6245
rect 4341 6205 4353 6239
rect 4387 6205 4399 6239
rect 4341 6199 4399 6205
rect 5169 6239 5227 6245
rect 5169 6205 5181 6239
rect 5215 6236 5227 6239
rect 5534 6236 5540 6248
rect 5215 6208 5540 6236
rect 5215 6205 5227 6208
rect 5169 6199 5227 6205
rect 3326 6128 3332 6180
rect 3384 6168 3390 6180
rect 3804 6168 3832 6199
rect 5534 6196 5540 6208
rect 5592 6196 5598 6248
rect 6104 6245 6132 6276
rect 6089 6239 6147 6245
rect 6089 6205 6101 6239
rect 6135 6205 6147 6239
rect 6089 6199 6147 6205
rect 6917 6239 6975 6245
rect 6917 6205 6929 6239
rect 6963 6236 6975 6239
rect 7006 6236 7012 6248
rect 6963 6208 7012 6236
rect 6963 6205 6975 6208
rect 6917 6199 6975 6205
rect 7006 6196 7012 6208
rect 7064 6196 7070 6248
rect 7101 6239 7159 6245
rect 7101 6205 7113 6239
rect 7147 6236 7159 6239
rect 7190 6236 7196 6248
rect 7147 6208 7196 6236
rect 7147 6205 7159 6208
rect 7101 6199 7159 6205
rect 7190 6196 7196 6208
rect 7248 6196 7254 6248
rect 7282 6196 7288 6248
rect 7340 6236 7346 6248
rect 7760 6245 7788 6276
rect 7852 6276 8616 6304
rect 7852 6248 7880 6276
rect 7619 6239 7677 6245
rect 7619 6236 7631 6239
rect 7340 6208 7631 6236
rect 7340 6196 7346 6208
rect 7619 6205 7631 6208
rect 7665 6205 7677 6239
rect 7619 6199 7677 6205
rect 7745 6239 7803 6245
rect 7745 6205 7757 6239
rect 7791 6205 7803 6239
rect 7745 6199 7803 6205
rect 7834 6196 7840 6248
rect 7892 6236 7898 6248
rect 8018 6236 8024 6248
rect 7892 6208 7937 6236
rect 7979 6208 8024 6236
rect 7892 6196 7898 6208
rect 8018 6196 8024 6208
rect 8076 6196 8082 6248
rect 8588 6245 8616 6276
rect 8573 6239 8631 6245
rect 8573 6205 8585 6239
rect 8619 6205 8631 6239
rect 8573 6199 8631 6205
rect 8662 6196 8668 6248
rect 8720 6236 8726 6248
rect 8956 6245 8984 6412
rect 10321 6409 10333 6412
rect 10367 6409 10379 6443
rect 10321 6403 10379 6409
rect 9033 6375 9091 6381
rect 9033 6341 9045 6375
rect 9079 6372 9091 6375
rect 9950 6372 9956 6384
rect 9079 6344 9956 6372
rect 9079 6341 9091 6344
rect 9033 6335 9091 6341
rect 9950 6332 9956 6344
rect 10008 6332 10014 6384
rect 11057 6375 11115 6381
rect 11057 6372 11069 6375
rect 10152 6344 11069 6372
rect 8849 6239 8907 6245
rect 8849 6236 8861 6239
rect 8720 6208 8861 6236
rect 8720 6196 8726 6208
rect 8849 6205 8861 6208
rect 8895 6205 8907 6239
rect 8849 6199 8907 6205
rect 8941 6239 8999 6245
rect 8941 6205 8953 6239
rect 8987 6205 8999 6239
rect 8941 6199 8999 6205
rect 5997 6171 6055 6177
rect 3384 6140 4844 6168
rect 3384 6128 3390 6140
rect 4816 6109 4844 6140
rect 5997 6137 6009 6171
rect 6043 6168 6055 6171
rect 8956 6168 8984 6199
rect 9122 6196 9128 6248
rect 9180 6236 9186 6248
rect 9723 6239 9781 6245
rect 9180 6208 9225 6236
rect 9180 6196 9186 6208
rect 9723 6205 9735 6239
rect 9769 6205 9781 6239
rect 9723 6199 9781 6205
rect 6043 6140 8984 6168
rect 6043 6137 6055 6140
rect 5997 6131 6055 6137
rect 7760 6112 7788 6140
rect 9030 6128 9036 6180
rect 9088 6168 9094 6180
rect 9738 6168 9766 6199
rect 9858 6196 9864 6248
rect 9916 6236 9922 6248
rect 10152 6245 10180 6344
rect 11057 6341 11069 6344
rect 11103 6341 11115 6375
rect 11057 6335 11115 6341
rect 10321 6307 10379 6313
rect 10321 6273 10333 6307
rect 10367 6304 10379 6307
rect 11977 6307 12035 6313
rect 10367 6276 10921 6304
rect 10367 6273 10379 6276
rect 10321 6267 10379 6273
rect 10137 6239 10195 6245
rect 10137 6236 10149 6239
rect 9916 6208 10149 6236
rect 9916 6196 9922 6208
rect 10137 6205 10149 6208
rect 10183 6205 10195 6239
rect 10502 6236 10508 6248
rect 10463 6208 10508 6236
rect 10137 6199 10195 6205
rect 10502 6196 10508 6208
rect 10560 6196 10566 6248
rect 10893 6245 10921 6276
rect 11977 6273 11989 6307
rect 12023 6304 12035 6307
rect 12710 6304 12716 6316
rect 12023 6276 12716 6304
rect 12023 6273 12035 6276
rect 11977 6267 12035 6273
rect 12710 6264 12716 6276
rect 12768 6304 12774 6316
rect 13262 6304 13268 6316
rect 12768 6276 13268 6304
rect 12768 6264 12774 6276
rect 13262 6264 13268 6276
rect 13320 6264 13326 6316
rect 10878 6239 10936 6245
rect 10878 6205 10890 6239
rect 10924 6205 10936 6239
rect 10878 6199 10936 6205
rect 12437 6239 12495 6245
rect 12437 6205 12449 6239
rect 12483 6236 12495 6239
rect 12894 6236 12900 6248
rect 12483 6208 12900 6236
rect 12483 6205 12495 6208
rect 12437 6199 12495 6205
rect 12894 6196 12900 6208
rect 12952 6236 12958 6248
rect 13357 6239 13415 6245
rect 13357 6236 13369 6239
rect 12952 6208 13369 6236
rect 12952 6196 12958 6208
rect 13357 6205 13369 6208
rect 13403 6205 13415 6239
rect 13357 6199 13415 6205
rect 10229 6171 10287 6177
rect 10229 6168 10241 6171
rect 9088 6140 10241 6168
rect 9088 6128 9094 6140
rect 10229 6137 10241 6140
rect 10275 6137 10287 6171
rect 10686 6168 10692 6180
rect 10647 6140 10692 6168
rect 10229 6131 10287 6137
rect 10686 6128 10692 6140
rect 10744 6128 10750 6180
rect 10778 6128 10784 6180
rect 10836 6168 10842 6180
rect 11793 6171 11851 6177
rect 11793 6168 11805 6171
rect 10836 6140 10881 6168
rect 10980 6140 11805 6168
rect 10836 6128 10842 6140
rect 4801 6103 4859 6109
rect 4801 6069 4813 6103
rect 4847 6069 4859 6103
rect 4801 6063 4859 6069
rect 7742 6060 7748 6112
rect 7800 6060 7806 6112
rect 9585 6103 9643 6109
rect 9585 6069 9597 6103
rect 9631 6100 9643 6103
rect 9858 6100 9864 6112
rect 9631 6072 9864 6100
rect 9631 6069 9643 6072
rect 9585 6063 9643 6069
rect 9858 6060 9864 6072
rect 9916 6060 9922 6112
rect 9950 6060 9956 6112
rect 10008 6100 10014 6112
rect 10980 6100 11008 6140
rect 11793 6137 11805 6140
rect 11839 6137 11851 6171
rect 11793 6131 11851 6137
rect 10008 6072 11008 6100
rect 10008 6060 10014 6072
rect 11146 6060 11152 6112
rect 11204 6100 11210 6112
rect 12253 6103 12311 6109
rect 12253 6100 12265 6103
rect 11204 6072 12265 6100
rect 11204 6060 11210 6072
rect 12253 6069 12265 6072
rect 12299 6069 12311 6103
rect 12253 6063 12311 6069
rect 12713 6103 12771 6109
rect 12713 6069 12725 6103
rect 12759 6100 12771 6103
rect 12802 6100 12808 6112
rect 12759 6072 12808 6100
rect 12759 6069 12771 6072
rect 12713 6063 12771 6069
rect 12802 6060 12808 6072
rect 12860 6060 12866 6112
rect 13170 6100 13176 6112
rect 13131 6072 13176 6100
rect 13170 6060 13176 6072
rect 13228 6060 13234 6112
rect 1104 6010 13892 6032
rect 1104 5958 8246 6010
rect 8298 5958 8310 6010
rect 8362 5958 8374 6010
rect 8426 5958 8438 6010
rect 8490 5958 13892 6010
rect 1104 5936 13892 5958
rect 1394 5896 1400 5908
rect 1355 5868 1400 5896
rect 1394 5856 1400 5868
rect 1452 5856 1458 5908
rect 1854 5896 1860 5908
rect 1815 5868 1860 5896
rect 1854 5856 1860 5868
rect 1912 5856 1918 5908
rect 5261 5899 5319 5905
rect 3160 5868 5212 5896
rect 2777 5831 2835 5837
rect 2777 5797 2789 5831
rect 2823 5828 2835 5831
rect 3050 5828 3056 5840
rect 2823 5800 3056 5828
rect 2823 5797 2835 5800
rect 2777 5791 2835 5797
rect 3050 5788 3056 5800
rect 3108 5788 3114 5840
rect 1765 5763 1823 5769
rect 1765 5729 1777 5763
rect 1811 5760 1823 5763
rect 3160 5760 3188 5868
rect 4617 5831 4675 5837
rect 4617 5797 4629 5831
rect 4663 5828 4675 5831
rect 4798 5828 4804 5840
rect 4663 5800 4804 5828
rect 4663 5797 4675 5800
rect 4617 5791 4675 5797
rect 4798 5788 4804 5800
rect 4856 5788 4862 5840
rect 5184 5828 5212 5868
rect 5261 5865 5273 5899
rect 5307 5896 5319 5899
rect 6730 5896 6736 5908
rect 5307 5868 6736 5896
rect 5307 5865 5319 5868
rect 5261 5859 5319 5865
rect 6730 5856 6736 5868
rect 6788 5896 6794 5908
rect 10778 5896 10784 5908
rect 6788 5868 8156 5896
rect 6788 5856 6794 5868
rect 6178 5828 6184 5840
rect 5184 5800 6184 5828
rect 6178 5788 6184 5800
rect 6236 5788 6242 5840
rect 6362 5788 6368 5840
rect 6420 5788 6426 5840
rect 7190 5788 7196 5840
rect 7248 5828 7254 5840
rect 7926 5828 7932 5840
rect 7248 5800 7932 5828
rect 7248 5788 7254 5800
rect 7926 5788 7932 5800
rect 7984 5788 7990 5840
rect 3326 5760 3332 5772
rect 1811 5732 3188 5760
rect 3287 5732 3332 5760
rect 1811 5729 1823 5732
rect 1765 5723 1823 5729
rect 3326 5720 3332 5732
rect 3384 5720 3390 5772
rect 3510 5720 3516 5772
rect 3568 5760 3574 5772
rect 4065 5763 4123 5769
rect 4065 5760 4077 5763
rect 3568 5732 4077 5760
rect 3568 5720 3574 5732
rect 4065 5729 4077 5732
rect 4111 5729 4123 5763
rect 4065 5723 4123 5729
rect 4525 5763 4583 5769
rect 4525 5729 4537 5763
rect 4571 5760 4583 5763
rect 4706 5760 4712 5772
rect 4571 5732 4712 5760
rect 4571 5729 4583 5732
rect 4525 5723 4583 5729
rect 4706 5720 4712 5732
rect 4764 5720 4770 5772
rect 5353 5763 5411 5769
rect 5353 5729 5365 5763
rect 5399 5729 5411 5763
rect 5626 5760 5632 5772
rect 5587 5732 5632 5760
rect 5353 5723 5411 5729
rect 2038 5692 2044 5704
rect 1999 5664 2044 5692
rect 2038 5652 2044 5664
rect 2096 5652 2102 5704
rect 2866 5692 2872 5704
rect 2827 5664 2872 5692
rect 2866 5652 2872 5664
rect 2924 5652 2930 5704
rect 5368 5692 5396 5723
rect 5626 5720 5632 5732
rect 5684 5720 5690 5772
rect 7834 5692 7840 5704
rect 5368 5664 7840 5692
rect 7834 5652 7840 5664
rect 7892 5652 7898 5704
rect 8128 5692 8156 5868
rect 9140 5868 10784 5896
rect 9030 5828 9036 5840
rect 8220 5800 9036 5828
rect 8220 5769 8248 5800
rect 9030 5788 9036 5800
rect 9088 5788 9094 5840
rect 8205 5763 8263 5769
rect 8205 5729 8217 5763
rect 8251 5729 8263 5763
rect 8205 5723 8263 5729
rect 8297 5763 8355 5769
rect 8297 5729 8309 5763
rect 8343 5729 8355 5763
rect 8297 5723 8355 5729
rect 8573 5763 8631 5769
rect 8573 5729 8585 5763
rect 8619 5760 8631 5763
rect 8754 5760 8760 5772
rect 8619 5732 8760 5760
rect 8619 5729 8631 5732
rect 8573 5723 8631 5729
rect 8312 5692 8340 5723
rect 8754 5720 8760 5732
rect 8812 5720 8818 5772
rect 9140 5769 9168 5868
rect 10778 5856 10784 5868
rect 10836 5856 10842 5908
rect 10962 5896 10968 5908
rect 10923 5868 10968 5896
rect 10962 5856 10968 5868
rect 11020 5856 11026 5908
rect 9217 5831 9275 5837
rect 9217 5797 9229 5831
rect 9263 5828 9275 5831
rect 9766 5828 9772 5840
rect 9263 5800 9772 5828
rect 9263 5797 9275 5800
rect 9217 5791 9275 5797
rect 9766 5788 9772 5800
rect 9824 5828 9830 5840
rect 10686 5828 10692 5840
rect 9824 5800 10692 5828
rect 9824 5788 9830 5800
rect 9125 5763 9183 5769
rect 9125 5729 9137 5763
rect 9171 5729 9183 5763
rect 9125 5723 9183 5729
rect 9493 5763 9551 5769
rect 9493 5729 9505 5763
rect 9539 5760 9551 5763
rect 9585 5763 9643 5769
rect 9585 5760 9597 5763
rect 9539 5732 9597 5760
rect 9539 5729 9551 5732
rect 9493 5723 9551 5729
rect 9585 5729 9597 5732
rect 9631 5729 9643 5763
rect 9858 5760 9864 5772
rect 9819 5732 9864 5760
rect 9585 5723 9643 5729
rect 8128 5664 8340 5692
rect 7852 5624 7880 5652
rect 8312 5624 8340 5664
rect 8662 5652 8668 5704
rect 8720 5692 8726 5704
rect 9140 5692 9168 5723
rect 9858 5720 9864 5732
rect 9916 5720 9922 5772
rect 10336 5769 10364 5800
rect 10686 5788 10692 5800
rect 10744 5788 10750 5840
rect 11057 5831 11115 5837
rect 11057 5797 11069 5831
rect 11103 5828 11115 5831
rect 11238 5828 11244 5840
rect 11103 5800 11244 5828
rect 11103 5797 11115 5800
rect 11057 5791 11115 5797
rect 11238 5788 11244 5800
rect 11296 5788 11302 5840
rect 11698 5828 11704 5840
rect 11659 5800 11704 5828
rect 11698 5788 11704 5800
rect 11756 5788 11762 5840
rect 13170 5828 13176 5840
rect 12926 5800 13176 5828
rect 13170 5788 13176 5800
rect 13228 5788 13234 5840
rect 10137 5763 10195 5769
rect 10137 5729 10149 5763
rect 10183 5729 10195 5763
rect 10137 5723 10195 5729
rect 10321 5763 10379 5769
rect 10321 5729 10333 5763
rect 10367 5729 10379 5763
rect 10321 5723 10379 5729
rect 8720 5664 9168 5692
rect 8720 5652 8726 5664
rect 9766 5652 9772 5704
rect 9824 5692 9830 5704
rect 9953 5695 10011 5701
rect 9953 5692 9965 5695
rect 9824 5664 9965 5692
rect 9824 5652 9830 5664
rect 9953 5661 9965 5664
rect 9999 5661 10011 5695
rect 9953 5655 10011 5661
rect 7852 5596 8156 5624
rect 8312 5596 8984 5624
rect 5534 5516 5540 5568
rect 5592 5556 5598 5568
rect 5886 5559 5944 5565
rect 5886 5556 5898 5559
rect 5592 5528 5898 5556
rect 5592 5516 5598 5528
rect 5886 5525 5898 5528
rect 5932 5525 5944 5559
rect 7374 5556 7380 5568
rect 7335 5528 7380 5556
rect 5886 5519 5944 5525
rect 7374 5516 7380 5528
rect 7432 5516 7438 5568
rect 8018 5556 8024 5568
rect 7979 5528 8024 5556
rect 8018 5516 8024 5528
rect 8076 5516 8082 5568
rect 8128 5556 8156 5596
rect 8478 5556 8484 5568
rect 8128 5528 8484 5556
rect 8478 5516 8484 5528
rect 8536 5516 8542 5568
rect 8956 5556 8984 5596
rect 9030 5584 9036 5636
rect 9088 5624 9094 5636
rect 9858 5624 9864 5636
rect 9088 5596 9864 5624
rect 9088 5584 9094 5596
rect 9858 5584 9864 5596
rect 9916 5584 9922 5636
rect 9493 5559 9551 5565
rect 9493 5556 9505 5559
rect 8956 5528 9505 5556
rect 9493 5525 9505 5528
rect 9539 5525 9551 5559
rect 9493 5519 9551 5525
rect 9582 5516 9588 5568
rect 9640 5556 9646 5568
rect 10152 5556 10180 5723
rect 10226 5652 10232 5704
rect 10284 5692 10290 5704
rect 11425 5695 11483 5701
rect 11425 5692 11437 5695
rect 10284 5664 11437 5692
rect 10284 5652 10290 5664
rect 11425 5661 11437 5664
rect 11471 5661 11483 5695
rect 11425 5655 11483 5661
rect 9640 5528 10180 5556
rect 11440 5556 11468 5655
rect 11514 5556 11520 5568
rect 11440 5528 11520 5556
rect 9640 5516 9646 5528
rect 11514 5516 11520 5528
rect 11572 5516 11578 5568
rect 13170 5556 13176 5568
rect 13131 5528 13176 5556
rect 13170 5516 13176 5528
rect 13228 5516 13234 5568
rect 1104 5466 13892 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 12246 5466
rect 12298 5414 12310 5466
rect 12362 5414 12374 5466
rect 12426 5414 12438 5466
rect 12490 5414 13892 5466
rect 1104 5392 13892 5414
rect 5626 5312 5632 5364
rect 5684 5352 5690 5364
rect 5994 5352 6000 5364
rect 5684 5324 6000 5352
rect 5684 5312 5690 5324
rect 5994 5312 6000 5324
rect 6052 5352 6058 5364
rect 7466 5352 7472 5364
rect 6052 5324 7472 5352
rect 6052 5312 6058 5324
rect 7466 5312 7472 5324
rect 7524 5352 7530 5364
rect 8754 5352 8760 5364
rect 7524 5324 8616 5352
rect 8715 5324 8760 5352
rect 7524 5312 7530 5324
rect 4338 5176 4344 5228
rect 4396 5216 4402 5228
rect 7285 5219 7343 5225
rect 4396 5188 6500 5216
rect 4396 5176 4402 5188
rect 1578 5148 1584 5160
rect 1539 5120 1584 5148
rect 1578 5108 1584 5120
rect 1636 5108 1642 5160
rect 3881 5151 3939 5157
rect 3881 5117 3893 5151
rect 3927 5148 3939 5151
rect 4062 5148 4068 5160
rect 3927 5120 4068 5148
rect 3927 5117 3939 5120
rect 3881 5111 3939 5117
rect 4062 5108 4068 5120
rect 4120 5108 4126 5160
rect 4614 5108 4620 5160
rect 4672 5108 4678 5160
rect 5994 5108 6000 5160
rect 6052 5148 6058 5160
rect 6472 5157 6500 5188
rect 7285 5185 7297 5219
rect 7331 5216 7343 5219
rect 8018 5216 8024 5228
rect 7331 5188 8024 5216
rect 7331 5185 7343 5188
rect 7285 5179 7343 5185
rect 8018 5176 8024 5188
rect 8076 5176 8082 5228
rect 8588 5216 8616 5324
rect 8754 5312 8760 5324
rect 8812 5312 8818 5364
rect 10226 5352 10232 5364
rect 9508 5324 10232 5352
rect 9398 5216 9404 5228
rect 8588 5188 9404 5216
rect 9398 5176 9404 5188
rect 9456 5216 9462 5228
rect 9508 5225 9536 5324
rect 10226 5312 10232 5324
rect 10284 5312 10290 5364
rect 10778 5312 10784 5364
rect 10836 5352 10842 5364
rect 11241 5355 11299 5361
rect 11241 5352 11253 5355
rect 10836 5324 11253 5352
rect 10836 5312 10842 5324
rect 11241 5321 11253 5324
rect 11287 5321 11299 5355
rect 11241 5315 11299 5321
rect 12529 5287 12587 5293
rect 12529 5284 12541 5287
rect 11900 5256 12541 5284
rect 9493 5219 9551 5225
rect 9493 5216 9505 5219
rect 9456 5188 9505 5216
rect 9456 5176 9462 5188
rect 9493 5185 9505 5188
rect 9539 5185 9551 5219
rect 9766 5216 9772 5228
rect 9727 5188 9772 5216
rect 9493 5179 9551 5185
rect 9766 5176 9772 5188
rect 9824 5176 9830 5228
rect 11900 5160 11928 5256
rect 12529 5253 12541 5256
rect 12575 5253 12587 5287
rect 12529 5247 12587 5253
rect 12434 5176 12440 5228
rect 12492 5216 12498 5228
rect 12693 5219 12751 5225
rect 12693 5216 12705 5219
rect 12492 5188 12705 5216
rect 12492 5176 12498 5188
rect 12693 5185 12705 5188
rect 12739 5216 12751 5219
rect 13170 5216 13176 5228
rect 12739 5188 13176 5216
rect 12739 5185 12751 5188
rect 12693 5179 12751 5185
rect 13170 5176 13176 5188
rect 13228 5176 13234 5228
rect 6457 5151 6515 5157
rect 6052 5120 6097 5148
rect 6052 5108 6058 5120
rect 6457 5117 6469 5151
rect 6503 5117 6515 5151
rect 11882 5148 11888 5160
rect 11843 5120 11888 5148
rect 6457 5111 6515 5117
rect 11882 5108 11888 5120
rect 11940 5108 11946 5160
rect 12805 5151 12863 5157
rect 12805 5117 12817 5151
rect 12851 5117 12863 5151
rect 12805 5111 12863 5117
rect 3602 5080 3608 5092
rect 1780 5052 2438 5080
rect 3563 5052 3608 5080
rect 1780 5021 1808 5052
rect 3602 5040 3608 5052
rect 3660 5040 3666 5092
rect 5718 5080 5724 5092
rect 5679 5052 5724 5080
rect 5718 5040 5724 5052
rect 5776 5040 5782 5092
rect 5810 5040 5816 5092
rect 5868 5080 5874 5092
rect 11146 5080 11152 5092
rect 5868 5052 7774 5080
rect 10994 5052 11152 5080
rect 5868 5040 5874 5052
rect 11146 5040 11152 5052
rect 11204 5040 11210 5092
rect 12820 5080 12848 5111
rect 13078 5080 13084 5092
rect 12820 5052 13084 5080
rect 13078 5040 13084 5052
rect 13136 5040 13142 5092
rect 1765 5015 1823 5021
rect 1765 4981 1777 5015
rect 1811 4981 1823 5015
rect 2130 5012 2136 5024
rect 2091 4984 2136 5012
rect 1765 4975 1823 4981
rect 2130 4972 2136 4984
rect 2188 4972 2194 5024
rect 4249 5015 4307 5021
rect 4249 4981 4261 5015
rect 4295 5012 4307 5015
rect 6362 5012 6368 5024
rect 4295 4984 6368 5012
rect 4295 4981 4307 4984
rect 4249 4975 4307 4981
rect 6362 4972 6368 4984
rect 6420 4972 6426 5024
rect 6546 5012 6552 5024
rect 6507 4984 6552 5012
rect 6546 4972 6552 4984
rect 6604 4972 6610 5024
rect 11790 5012 11796 5024
rect 11751 4984 11796 5012
rect 11790 4972 11796 4984
rect 11848 4972 11854 5024
rect 1104 4922 13892 4944
rect 1104 4870 8246 4922
rect 8298 4870 8310 4922
rect 8362 4870 8374 4922
rect 8426 4870 8438 4922
rect 8490 4870 13892 4922
rect 1104 4848 13892 4870
rect 2424 4780 3556 4808
rect 1581 4675 1639 4681
rect 1581 4641 1593 4675
rect 1627 4641 1639 4675
rect 2038 4672 2044 4684
rect 1999 4644 2044 4672
rect 1581 4635 1639 4641
rect 1596 4604 1624 4635
rect 2038 4632 2044 4644
rect 2096 4632 2102 4684
rect 2130 4632 2136 4684
rect 2188 4672 2194 4684
rect 2424 4681 2452 4780
rect 3528 4740 3556 4780
rect 3602 4768 3608 4820
rect 3660 4808 3666 4820
rect 3956 4811 4014 4817
rect 3956 4808 3968 4811
rect 3660 4780 3968 4808
rect 3660 4768 3666 4780
rect 3956 4777 3968 4780
rect 4002 4777 4014 4811
rect 3956 4771 4014 4777
rect 4154 4768 4160 4820
rect 4212 4808 4218 4820
rect 5261 4811 5319 4817
rect 4212 4780 5212 4808
rect 4212 4768 4218 4780
rect 4249 4743 4307 4749
rect 4249 4740 4261 4743
rect 3528 4712 4261 4740
rect 2409 4675 2467 4681
rect 2409 4672 2421 4675
rect 2188 4644 2421 4672
rect 2188 4632 2194 4644
rect 2409 4641 2421 4644
rect 2455 4641 2467 4675
rect 2409 4635 2467 4641
rect 2685 4675 2743 4681
rect 2685 4641 2697 4675
rect 2731 4672 2743 4675
rect 3329 4675 3387 4681
rect 3329 4672 3341 4675
rect 2731 4644 3341 4672
rect 2731 4641 2743 4644
rect 2685 4635 2743 4641
rect 3329 4641 3341 4644
rect 3375 4641 3387 4675
rect 3329 4635 3387 4641
rect 1946 4604 1952 4616
rect 1596 4576 1952 4604
rect 1946 4564 1952 4576
rect 2004 4564 2010 4616
rect 2317 4607 2375 4613
rect 2317 4573 2329 4607
rect 2363 4604 2375 4607
rect 2958 4604 2964 4616
rect 2363 4576 2964 4604
rect 2363 4573 2375 4576
rect 2317 4567 2375 4573
rect 2958 4564 2964 4576
rect 3016 4564 3022 4616
rect 3344 4604 3372 4635
rect 3418 4632 3424 4684
rect 3476 4672 3482 4684
rect 3528 4681 3556 4712
rect 4249 4709 4261 4712
rect 4295 4709 4307 4743
rect 5184 4740 5212 4780
rect 5261 4777 5273 4811
rect 5307 4808 5319 4811
rect 5718 4808 5724 4820
rect 5307 4780 5724 4808
rect 5307 4777 5319 4780
rect 5261 4771 5319 4777
rect 5718 4768 5724 4780
rect 5776 4768 5782 4820
rect 5813 4811 5871 4817
rect 5813 4777 5825 4811
rect 5859 4808 5871 4811
rect 6641 4811 6699 4817
rect 6641 4808 6653 4811
rect 5859 4780 6653 4808
rect 5859 4777 5871 4780
rect 5813 4771 5871 4777
rect 6641 4777 6653 4780
rect 6687 4777 6699 4811
rect 8846 4808 8852 4820
rect 6641 4771 6699 4777
rect 8312 4780 8852 4808
rect 5350 4740 5356 4752
rect 5184 4712 5356 4740
rect 4249 4703 4307 4709
rect 5350 4700 5356 4712
rect 5408 4740 5414 4752
rect 6273 4743 6331 4749
rect 5408 4712 6172 4740
rect 5408 4700 5414 4712
rect 4154 4681 4160 4684
rect 3513 4675 3571 4681
rect 3513 4672 3525 4675
rect 3476 4644 3525 4672
rect 3476 4632 3482 4644
rect 3513 4641 3525 4644
rect 3559 4641 3571 4675
rect 3513 4635 3571 4641
rect 4152 4635 4160 4681
rect 4212 4672 4218 4684
rect 4338 4672 4344 4684
rect 4212 4644 4252 4672
rect 4299 4644 4344 4672
rect 4154 4632 4160 4635
rect 4212 4632 4218 4644
rect 4338 4632 4344 4644
rect 4396 4632 4402 4684
rect 6144 4681 6172 4712
rect 6273 4709 6285 4743
rect 6319 4740 6331 4743
rect 6730 4740 6736 4752
rect 6319 4712 6736 4740
rect 6319 4709 6331 4712
rect 6273 4703 6331 4709
rect 6730 4700 6736 4712
rect 6788 4740 6794 4752
rect 6788 4712 7328 4740
rect 6788 4700 6794 4712
rect 4525 4675 4583 4681
rect 4525 4641 4537 4675
rect 4571 4672 4583 4675
rect 4985 4675 5043 4681
rect 4571 4644 4752 4672
rect 4571 4641 4583 4644
rect 4525 4635 4583 4641
rect 3878 4604 3884 4616
rect 3344 4576 3884 4604
rect 3878 4564 3884 4576
rect 3936 4604 3942 4616
rect 4356 4604 4384 4632
rect 3936 4576 4384 4604
rect 3936 4564 3942 4576
rect 1489 4539 1547 4545
rect 1489 4505 1501 4539
rect 1535 4536 1547 4539
rect 3053 4539 3111 4545
rect 1535 4508 3004 4536
rect 1535 4505 1547 4508
rect 1489 4499 1547 4505
rect 1949 4471 2007 4477
rect 1949 4437 1961 4471
rect 1995 4468 2007 4471
rect 2866 4468 2872 4480
rect 1995 4440 2872 4468
rect 1995 4437 2007 4440
rect 1949 4431 2007 4437
rect 2866 4428 2872 4440
rect 2924 4428 2930 4480
rect 2976 4468 3004 4508
rect 3053 4505 3065 4539
rect 3099 4536 3111 4539
rect 4614 4536 4620 4548
rect 3099 4508 4620 4536
rect 3099 4505 3111 4508
rect 3053 4499 3111 4505
rect 4614 4496 4620 4508
rect 4672 4496 4678 4548
rect 4724 4536 4752 4644
rect 4985 4641 4997 4675
rect 5031 4672 5043 4675
rect 6129 4675 6187 4681
rect 5031 4644 6040 4672
rect 5031 4641 5043 4644
rect 4985 4635 5043 4641
rect 4801 4607 4859 4613
rect 4801 4573 4813 4607
rect 4847 4604 4859 4607
rect 4890 4604 4896 4616
rect 4847 4576 4896 4604
rect 4847 4573 4859 4576
rect 4801 4567 4859 4573
rect 4890 4564 4896 4576
rect 4948 4564 4954 4616
rect 5353 4607 5411 4613
rect 5353 4573 5365 4607
rect 5399 4604 5411 4607
rect 5718 4604 5724 4616
rect 5399 4576 5724 4604
rect 5399 4573 5411 4576
rect 5353 4567 5411 4573
rect 5368 4536 5396 4567
rect 5718 4564 5724 4576
rect 5776 4604 5782 4616
rect 5813 4607 5871 4613
rect 5813 4604 5825 4607
rect 5776 4576 5825 4604
rect 5776 4564 5782 4576
rect 5813 4573 5825 4576
rect 5859 4573 5871 4607
rect 6012 4604 6040 4644
rect 6129 4641 6141 4675
rect 6175 4641 6187 4675
rect 6362 4672 6368 4684
rect 6323 4644 6368 4672
rect 6129 4635 6187 4641
rect 6362 4632 6368 4644
rect 6420 4632 6426 4684
rect 6549 4675 6607 4681
rect 6549 4641 6561 4675
rect 6595 4672 6607 4675
rect 6641 4675 6699 4681
rect 6641 4672 6653 4675
rect 6595 4644 6653 4672
rect 6595 4641 6607 4644
rect 6549 4635 6607 4641
rect 6641 4641 6653 4644
rect 6687 4641 6699 4675
rect 6822 4672 6828 4684
rect 6783 4644 6828 4672
rect 6641 4635 6699 4641
rect 6822 4632 6828 4644
rect 6880 4632 6886 4684
rect 7300 4681 7328 4712
rect 7285 4675 7343 4681
rect 7285 4641 7297 4675
rect 7331 4672 7343 4675
rect 7374 4672 7380 4684
rect 7331 4644 7380 4672
rect 7331 4641 7343 4644
rect 7285 4635 7343 4641
rect 7374 4632 7380 4644
rect 7432 4632 7438 4684
rect 7650 4632 7656 4684
rect 7708 4672 7714 4684
rect 8312 4681 8340 4780
rect 8846 4768 8852 4780
rect 8904 4768 8910 4820
rect 13078 4768 13084 4820
rect 13136 4808 13142 4820
rect 13265 4811 13323 4817
rect 13265 4808 13277 4811
rect 13136 4780 13277 4808
rect 13136 4768 13142 4780
rect 13265 4777 13277 4780
rect 13311 4777 13323 4811
rect 13265 4771 13323 4777
rect 9122 4740 9128 4752
rect 9083 4712 9128 4740
rect 9122 4700 9128 4712
rect 9180 4700 9186 4752
rect 12802 4700 12808 4752
rect 12860 4700 12866 4752
rect 8021 4675 8079 4681
rect 8021 4672 8033 4675
rect 7708 4644 8033 4672
rect 7708 4632 7714 4644
rect 8021 4641 8033 4644
rect 8067 4641 8079 4675
rect 8021 4635 8079 4641
rect 8297 4675 8355 4681
rect 8297 4641 8309 4675
rect 8343 4641 8355 4675
rect 8297 4635 8355 4641
rect 8481 4675 8539 4681
rect 8481 4641 8493 4675
rect 8527 4672 8539 4675
rect 8662 4672 8668 4684
rect 8527 4644 8668 4672
rect 8527 4641 8539 4644
rect 8481 4635 8539 4641
rect 8662 4632 8668 4644
rect 8720 4632 8726 4684
rect 8846 4632 8852 4684
rect 8904 4672 8910 4684
rect 9309 4675 9367 4681
rect 9309 4672 9321 4675
rect 8904 4644 9321 4672
rect 8904 4632 8910 4644
rect 9309 4641 9321 4644
rect 9355 4641 9367 4675
rect 9309 4635 9367 4641
rect 9678 4675 9736 4681
rect 9678 4641 9690 4675
rect 9724 4641 9736 4675
rect 9858 4672 9864 4684
rect 9819 4644 9864 4672
rect 9678 4635 9736 4641
rect 6917 4607 6975 4613
rect 6917 4604 6929 4607
rect 6012 4576 6929 4604
rect 5813 4567 5871 4573
rect 6917 4573 6929 4576
rect 6963 4604 6975 4607
rect 7006 4604 7012 4616
rect 6963 4576 7012 4604
rect 6963 4573 6975 4576
rect 6917 4567 6975 4573
rect 7006 4564 7012 4576
rect 7064 4564 7070 4616
rect 8754 4604 8760 4616
rect 8496 4576 8760 4604
rect 4724 4508 5396 4536
rect 5534 4496 5540 4548
rect 5592 4536 5598 4548
rect 5997 4539 6055 4545
rect 5997 4536 6009 4539
rect 5592 4508 6009 4536
rect 5592 4496 5598 4508
rect 5997 4505 6009 4508
rect 6043 4505 6055 4539
rect 7929 4539 7987 4545
rect 5997 4499 6055 4505
rect 6840 4508 7880 4536
rect 6840 4468 6868 4508
rect 7374 4468 7380 4480
rect 2976 4440 6868 4468
rect 7335 4440 7380 4468
rect 7374 4428 7380 4440
rect 7432 4428 7438 4480
rect 7852 4468 7880 4508
rect 7929 4505 7941 4539
rect 7975 4536 7987 4539
rect 7975 4508 8432 4536
rect 7975 4505 7987 4508
rect 7929 4499 7987 4505
rect 8404 4480 8432 4508
rect 8110 4468 8116 4480
rect 7852 4440 8116 4468
rect 8110 4428 8116 4440
rect 8168 4428 8174 4480
rect 8386 4428 8392 4480
rect 8444 4428 8450 4480
rect 8496 4477 8524 4576
rect 8754 4564 8760 4576
rect 8812 4564 8818 4616
rect 9490 4604 9496 4616
rect 9451 4576 9496 4604
rect 9490 4564 9496 4576
rect 9548 4564 9554 4616
rect 9585 4607 9643 4613
rect 9585 4573 9597 4607
rect 9631 4573 9643 4607
rect 9585 4567 9643 4573
rect 8665 4539 8723 4545
rect 8665 4505 8677 4539
rect 8711 4536 8723 4539
rect 9600 4536 9628 4567
rect 8711 4508 9628 4536
rect 9693 4536 9721 4635
rect 9858 4632 9864 4644
rect 9916 4632 9922 4684
rect 10505 4675 10563 4681
rect 10505 4641 10517 4675
rect 10551 4672 10563 4675
rect 10594 4672 10600 4684
rect 10551 4644 10600 4672
rect 10551 4641 10563 4644
rect 10505 4635 10563 4641
rect 10594 4632 10600 4644
rect 10652 4632 10658 4684
rect 10965 4675 11023 4681
rect 10965 4641 10977 4675
rect 11011 4672 11023 4675
rect 11054 4672 11060 4684
rect 11011 4644 11060 4672
rect 11011 4641 11023 4644
rect 10965 4635 11023 4641
rect 11054 4632 11060 4644
rect 11112 4632 11118 4684
rect 11514 4672 11520 4684
rect 11475 4644 11520 4672
rect 11514 4632 11520 4644
rect 11572 4632 11578 4684
rect 10134 4604 10140 4616
rect 10095 4576 10140 4604
rect 10134 4564 10140 4576
rect 10192 4564 10198 4616
rect 10686 4604 10692 4616
rect 10647 4576 10692 4604
rect 10686 4564 10692 4576
rect 10744 4564 10750 4616
rect 11793 4607 11851 4613
rect 11793 4573 11805 4607
rect 11839 4604 11851 4607
rect 12434 4604 12440 4616
rect 11839 4576 12440 4604
rect 11839 4573 11851 4576
rect 11793 4567 11851 4573
rect 12434 4564 12440 4576
rect 12492 4564 12498 4616
rect 9766 4536 9772 4548
rect 9693 4508 9772 4536
rect 8711 4505 8723 4508
rect 8665 4499 8723 4505
rect 9766 4496 9772 4508
rect 9824 4536 9830 4548
rect 10042 4536 10048 4548
rect 9824 4508 10048 4536
rect 9824 4496 9830 4508
rect 10042 4496 10048 4508
rect 10100 4496 10106 4548
rect 10229 4539 10287 4545
rect 10229 4505 10241 4539
rect 10275 4505 10287 4539
rect 10229 4499 10287 4505
rect 8481 4471 8539 4477
rect 8481 4437 8493 4471
rect 8527 4437 8539 4471
rect 8481 4431 8539 4437
rect 8754 4428 8760 4480
rect 8812 4468 8818 4480
rect 10244 4468 10272 4499
rect 11054 4468 11060 4480
rect 8812 4440 10272 4468
rect 11015 4440 11060 4468
rect 8812 4428 8818 4440
rect 11054 4428 11060 4440
rect 11112 4428 11118 4480
rect 1104 4378 13892 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 12246 4378
rect 12298 4326 12310 4378
rect 12362 4326 12374 4378
rect 12426 4326 12438 4378
rect 12490 4326 13892 4378
rect 1104 4304 13892 4326
rect 2866 4224 2872 4276
rect 2924 4264 2930 4276
rect 3053 4267 3111 4273
rect 3053 4264 3065 4267
rect 2924 4236 3065 4264
rect 2924 4224 2930 4236
rect 3053 4233 3065 4236
rect 3099 4233 3111 4267
rect 9756 4267 9814 4273
rect 3053 4227 3111 4233
rect 4080 4236 4476 4264
rect 2038 4156 2044 4208
rect 2096 4196 2102 4208
rect 4080 4196 4108 4236
rect 4448 4208 4476 4236
rect 9756 4233 9768 4267
rect 9802 4264 9814 4267
rect 11793 4267 11851 4273
rect 11793 4264 11805 4267
rect 9802 4236 11805 4264
rect 9802 4233 9814 4236
rect 9756 4227 9814 4233
rect 11793 4233 11805 4236
rect 11839 4233 11851 4267
rect 11793 4227 11851 4233
rect 2096 4168 4108 4196
rect 2096 4156 2102 4168
rect 4430 4156 4436 4208
rect 4488 4156 4494 4208
rect 11882 4156 11888 4208
rect 11940 4196 11946 4208
rect 11940 4168 12296 4196
rect 11940 4156 11946 4168
rect 474 4088 480 4140
rect 532 4128 538 4140
rect 1486 4128 1492 4140
rect 532 4100 1492 4128
rect 532 4088 538 4100
rect 1486 4088 1492 4100
rect 1544 4088 1550 4140
rect 8110 4128 8116 4140
rect 1780 4100 7972 4128
rect 8071 4100 8116 4128
rect 1780 4072 1808 4100
rect 1762 4060 1768 4072
rect 1675 4032 1768 4060
rect 1762 4020 1768 4032
rect 1820 4020 1826 4072
rect 1946 4060 1952 4072
rect 1907 4032 1952 4060
rect 1946 4020 1952 4032
rect 2004 4020 2010 4072
rect 2041 4063 2099 4069
rect 2041 4029 2053 4063
rect 2087 4029 2099 4063
rect 2041 4023 2099 4029
rect 2056 3924 2084 4023
rect 2130 4020 2136 4072
rect 2188 4060 2194 4072
rect 2958 4060 2964 4072
rect 2188 4032 2233 4060
rect 2919 4032 2964 4060
rect 2188 4020 2194 4032
rect 2958 4020 2964 4032
rect 3016 4020 3022 4072
rect 3483 4063 3541 4069
rect 3483 4029 3495 4063
rect 3529 4060 3541 4063
rect 3878 4060 3884 4072
rect 3529 4032 3884 4060
rect 3529 4029 3541 4032
rect 3483 4023 3541 4029
rect 3878 4020 3884 4032
rect 3936 4020 3942 4072
rect 5905 4063 5963 4069
rect 5905 4029 5917 4063
rect 5951 4060 5963 4063
rect 5994 4060 6000 4072
rect 5951 4032 6000 4060
rect 5951 4029 5963 4032
rect 5905 4023 5963 4029
rect 5994 4020 6000 4032
rect 6052 4020 6058 4072
rect 6730 4069 6736 4072
rect 6728 4060 6736 4069
rect 6691 4032 6736 4060
rect 6728 4023 6736 4032
rect 6730 4020 6736 4023
rect 6788 4020 6794 4072
rect 7098 4060 7104 4072
rect 7011 4032 7104 4060
rect 7098 4020 7104 4032
rect 7156 4060 7162 4072
rect 7374 4060 7380 4072
rect 7156 4032 7380 4060
rect 7156 4020 7162 4032
rect 7374 4020 7380 4032
rect 7432 4020 7438 4072
rect 7944 4069 7972 4100
rect 8110 4088 8116 4100
rect 8168 4088 8174 4140
rect 8205 4131 8263 4137
rect 8205 4097 8217 4131
rect 8251 4128 8263 4131
rect 8754 4128 8760 4140
rect 8251 4100 8760 4128
rect 8251 4097 8263 4100
rect 8205 4091 8263 4097
rect 8754 4088 8760 4100
rect 8812 4088 8818 4140
rect 9125 4131 9183 4137
rect 9125 4097 9137 4131
rect 9171 4128 9183 4131
rect 9766 4128 9772 4140
rect 9171 4100 9772 4128
rect 9171 4097 9183 4100
rect 9125 4091 9183 4097
rect 9766 4088 9772 4100
rect 9824 4088 9830 4140
rect 11238 4128 11244 4140
rect 11151 4100 11244 4128
rect 11238 4088 11244 4100
rect 11296 4128 11302 4140
rect 11296 4100 12204 4128
rect 11296 4088 11302 4100
rect 8386 4069 8392 4072
rect 7929 4063 7987 4069
rect 7929 4029 7941 4063
rect 7975 4029 7987 4063
rect 7929 4023 7987 4029
rect 8333 4063 8392 4069
rect 8333 4029 8345 4063
rect 8379 4029 8392 4063
rect 8333 4023 8392 4029
rect 8386 4020 8392 4023
rect 8444 4020 8450 4072
rect 8481 4063 8539 4069
rect 8481 4029 8493 4063
rect 8527 4060 8539 4063
rect 8570 4060 8576 4072
rect 8527 4032 8576 4060
rect 8527 4029 8539 4032
rect 8481 4023 8539 4029
rect 8570 4020 8576 4032
rect 8628 4020 8634 4072
rect 9398 4020 9404 4072
rect 9456 4060 9462 4072
rect 9493 4063 9551 4069
rect 9493 4060 9505 4063
rect 9456 4032 9505 4060
rect 9456 4020 9462 4032
rect 9493 4029 9505 4032
rect 9539 4029 9551 4063
rect 9493 4023 9551 4029
rect 11790 4020 11796 4072
rect 11848 4060 11854 4072
rect 12176 4069 12204 4100
rect 11925 4063 11983 4069
rect 11925 4060 11937 4063
rect 11848 4032 11937 4060
rect 11848 4020 11854 4032
rect 11925 4029 11937 4032
rect 11971 4029 11983 4063
rect 11925 4023 11983 4029
rect 12161 4063 12219 4069
rect 12161 4029 12173 4063
rect 12207 4029 12219 4063
rect 12268 4060 12296 4168
rect 12894 4156 12900 4208
rect 12952 4156 12958 4208
rect 12912 4128 12940 4156
rect 12912 4100 13124 4128
rect 13096 4072 13124 4100
rect 12345 4063 12403 4069
rect 12345 4060 12357 4063
rect 12268 4032 12357 4060
rect 12161 4023 12219 4029
rect 12345 4029 12357 4032
rect 12391 4029 12403 4063
rect 12345 4023 12403 4029
rect 12621 4063 12679 4069
rect 12621 4029 12633 4063
rect 12667 4060 12679 4063
rect 12894 4060 12900 4072
rect 12667 4032 12900 4060
rect 12667 4029 12679 4032
rect 12621 4023 12679 4029
rect 12894 4020 12900 4032
rect 12952 4020 12958 4072
rect 13078 4020 13084 4072
rect 13136 4060 13142 4072
rect 13265 4063 13323 4069
rect 13265 4060 13277 4063
rect 13136 4032 13277 4060
rect 13136 4020 13142 4032
rect 13265 4029 13277 4032
rect 13311 4029 13323 4063
rect 13265 4023 13323 4029
rect 2409 3995 2467 4001
rect 2409 3961 2421 3995
rect 2455 3992 2467 3995
rect 3326 3992 3332 4004
rect 2455 3964 3332 3992
rect 2455 3961 2467 3964
rect 2409 3955 2467 3961
rect 3326 3952 3332 3964
rect 3384 3952 3390 4004
rect 5626 3992 5632 4004
rect 3620 3964 4292 3992
rect 2222 3924 2228 3936
rect 2056 3896 2228 3924
rect 2222 3884 2228 3896
rect 2280 3884 2286 3936
rect 3418 3924 3424 3936
rect 3379 3896 3424 3924
rect 3418 3884 3424 3896
rect 3476 3924 3482 3936
rect 3620 3933 3648 3964
rect 3605 3927 3663 3933
rect 3605 3924 3617 3927
rect 3476 3896 3617 3924
rect 3476 3884 3482 3896
rect 3605 3893 3617 3896
rect 3651 3893 3663 3927
rect 3605 3887 3663 3893
rect 3878 3884 3884 3936
rect 3936 3924 3942 3936
rect 4157 3927 4215 3933
rect 4157 3924 4169 3927
rect 3936 3896 4169 3924
rect 3936 3884 3942 3896
rect 4157 3893 4169 3896
rect 4203 3893 4215 3927
rect 4264 3924 4292 3964
rect 4724 3936 4752 3978
rect 5587 3964 5632 3992
rect 5626 3952 5632 3964
rect 5684 3952 5690 4004
rect 6362 3952 6368 4004
rect 6420 3992 6426 4004
rect 6822 3992 6828 4004
rect 6420 3964 6828 3992
rect 6420 3952 6426 3964
rect 6822 3952 6828 3964
rect 6880 3952 6886 4004
rect 6917 3995 6975 4001
rect 6917 3961 6929 3995
rect 6963 3992 6975 3995
rect 7006 3992 7012 4004
rect 6963 3964 7012 3992
rect 6963 3961 6975 3964
rect 6917 3955 6975 3961
rect 7006 3952 7012 3964
rect 7064 3952 7070 4004
rect 8754 3992 8760 4004
rect 8715 3964 8760 3992
rect 8754 3952 8760 3964
rect 8812 3952 8818 4004
rect 8941 3995 8999 4001
rect 8941 3961 8953 3995
rect 8987 3961 8999 3995
rect 12066 3992 12072 4004
rect 10994 3964 11376 3992
rect 12027 3964 12072 3992
rect 8941 3955 8999 3961
rect 4614 3924 4620 3936
rect 4264 3896 4620 3924
rect 4157 3887 4215 3893
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 4706 3884 4712 3936
rect 4764 3884 4770 3936
rect 4982 3884 4988 3936
rect 5040 3924 5046 3936
rect 6270 3924 6276 3936
rect 5040 3896 6276 3924
rect 5040 3884 5046 3896
rect 6270 3884 6276 3896
rect 6328 3884 6334 3936
rect 6541 3927 6599 3933
rect 6541 3893 6553 3927
rect 6587 3924 6599 3927
rect 6730 3924 6736 3936
rect 6587 3896 6736 3924
rect 6587 3893 6599 3896
rect 6541 3887 6599 3893
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 7837 3927 7895 3933
rect 7837 3893 7849 3927
rect 7883 3924 7895 3927
rect 8956 3924 8984 3955
rect 7883 3896 8984 3924
rect 11348 3924 11376 3964
rect 12066 3952 12072 3964
rect 12124 3952 12130 4004
rect 12406 3964 13124 3992
rect 12406 3924 12434 3964
rect 12710 3924 12716 3936
rect 11348 3896 12434 3924
rect 12671 3896 12716 3924
rect 7883 3893 7895 3896
rect 7837 3887 7895 3893
rect 12710 3884 12716 3896
rect 12768 3884 12774 3936
rect 13096 3933 13124 3964
rect 13081 3927 13139 3933
rect 13081 3893 13093 3927
rect 13127 3893 13139 3927
rect 13081 3887 13139 3893
rect 1104 3834 13892 3856
rect 1104 3782 8246 3834
rect 8298 3782 8310 3834
rect 8362 3782 8374 3834
rect 8426 3782 8438 3834
rect 8490 3782 13892 3834
rect 1104 3760 13892 3782
rect 2593 3723 2651 3729
rect 2593 3689 2605 3723
rect 2639 3689 2651 3723
rect 5350 3720 5356 3732
rect 5311 3692 5356 3720
rect 2593 3683 2651 3689
rect 2608 3652 2636 3683
rect 5350 3680 5356 3692
rect 5408 3680 5414 3732
rect 5442 3680 5448 3732
rect 5500 3720 5506 3732
rect 5626 3720 5632 3732
rect 5500 3692 5545 3720
rect 5587 3692 5632 3720
rect 5500 3680 5506 3692
rect 5626 3680 5632 3692
rect 5684 3680 5690 3732
rect 9122 3720 9128 3732
rect 5736 3692 9128 3720
rect 3145 3655 3203 3661
rect 3145 3652 3157 3655
rect 1504 3624 2636 3652
rect 2884 3624 3157 3652
rect 1504 3596 1532 3624
rect 1486 3584 1492 3596
rect 1399 3556 1492 3584
rect 1486 3544 1492 3556
rect 1544 3544 1550 3596
rect 1670 3584 1676 3596
rect 1631 3556 1676 3584
rect 1670 3544 1676 3556
rect 1728 3544 1734 3596
rect 1854 3544 1860 3596
rect 1912 3584 1918 3596
rect 1949 3587 2007 3593
rect 1949 3584 1961 3587
rect 1912 3556 1961 3584
rect 1912 3544 1918 3556
rect 1949 3553 1961 3556
rect 1995 3584 2007 3587
rect 2038 3584 2044 3596
rect 1995 3556 2044 3584
rect 1995 3553 2007 3556
rect 1949 3547 2007 3553
rect 2038 3544 2044 3556
rect 2096 3544 2102 3596
rect 2222 3584 2228 3596
rect 2135 3556 2228 3584
rect 2222 3544 2228 3556
rect 2280 3544 2286 3596
rect 2884 3593 2912 3624
rect 3145 3621 3157 3624
rect 3191 3652 3203 3655
rect 4614 3652 4620 3664
rect 3191 3624 4620 3652
rect 3191 3621 3203 3624
rect 3145 3615 3203 3621
rect 4614 3612 4620 3624
rect 4672 3612 4678 3664
rect 5736 3652 5764 3692
rect 9122 3680 9128 3692
rect 9180 3680 9186 3732
rect 10134 3720 10140 3732
rect 9692 3692 10140 3720
rect 7006 3652 7012 3664
rect 5092 3624 5764 3652
rect 6932 3624 7012 3652
rect 2869 3587 2927 3593
rect 2869 3553 2881 3587
rect 2915 3553 2927 3587
rect 2869 3547 2927 3553
rect 3050 3544 3056 3596
rect 3108 3584 3114 3596
rect 3237 3587 3295 3593
rect 3237 3584 3249 3587
rect 3108 3556 3249 3584
rect 3108 3544 3114 3556
rect 3237 3553 3249 3556
rect 3283 3553 3295 3587
rect 3237 3547 3295 3553
rect 4249 3587 4307 3593
rect 4249 3553 4261 3587
rect 4295 3584 4307 3587
rect 4522 3584 4528 3596
rect 4295 3556 4528 3584
rect 4295 3553 4307 3556
rect 4249 3547 4307 3553
rect 4522 3544 4528 3556
rect 4580 3544 4586 3596
rect 1762 3408 1768 3460
rect 1820 3448 1826 3460
rect 1857 3451 1915 3457
rect 1857 3448 1869 3451
rect 1820 3420 1869 3448
rect 1820 3408 1826 3420
rect 1857 3417 1869 3420
rect 1903 3417 1915 3451
rect 2240 3448 2268 3544
rect 2757 3519 2815 3525
rect 2757 3485 2769 3519
rect 2803 3516 2815 3519
rect 3068 3516 3096 3544
rect 2803 3488 3096 3516
rect 2803 3485 2815 3488
rect 2757 3479 2815 3485
rect 3326 3476 3332 3528
rect 3384 3516 3390 3528
rect 4137 3519 4195 3525
rect 3384 3488 4108 3516
rect 3384 3476 3390 3488
rect 3973 3451 4031 3457
rect 3973 3448 3985 3451
rect 2240 3420 3985 3448
rect 1857 3411 1915 3417
rect 3973 3417 3985 3420
rect 4019 3417 4031 3451
rect 4080 3448 4108 3488
rect 4137 3485 4149 3519
rect 4183 3516 4195 3519
rect 4430 3516 4436 3528
rect 4183 3488 4436 3516
rect 4183 3485 4195 3488
rect 4137 3479 4195 3485
rect 4430 3476 4436 3488
rect 4488 3516 4494 3528
rect 4617 3519 4675 3525
rect 4617 3516 4629 3519
rect 4488 3488 4629 3516
rect 4488 3476 4494 3488
rect 4617 3485 4629 3488
rect 4663 3516 4675 3519
rect 5092 3516 5120 3624
rect 5169 3587 5227 3593
rect 5169 3553 5181 3587
rect 5215 3553 5227 3587
rect 5534 3584 5540 3596
rect 5495 3556 5540 3584
rect 5169 3547 5227 3553
rect 4663 3488 5120 3516
rect 5184 3516 5212 3547
rect 5534 3544 5540 3556
rect 5592 3544 5598 3596
rect 5902 3544 5908 3596
rect 5960 3584 5966 3596
rect 6273 3587 6331 3593
rect 6273 3584 6285 3587
rect 5960 3556 6285 3584
rect 5960 3544 5966 3556
rect 6273 3553 6285 3556
rect 6319 3553 6331 3587
rect 6273 3547 6331 3553
rect 6457 3587 6515 3593
rect 6457 3553 6469 3587
rect 6503 3584 6515 3587
rect 6546 3584 6552 3596
rect 6503 3556 6552 3584
rect 6503 3553 6515 3556
rect 6457 3547 6515 3553
rect 6546 3544 6552 3556
rect 6604 3544 6610 3596
rect 6932 3593 6960 3624
rect 7006 3612 7012 3624
rect 7064 3612 7070 3664
rect 7484 3624 8248 3652
rect 7484 3596 7512 3624
rect 6917 3587 6975 3593
rect 6917 3553 6929 3587
rect 6963 3553 6975 3587
rect 7098 3584 7104 3596
rect 7059 3556 7104 3584
rect 6917 3547 6975 3553
rect 7098 3544 7104 3556
rect 7156 3544 7162 3596
rect 7466 3584 7472 3596
rect 7427 3556 7472 3584
rect 7466 3544 7472 3556
rect 7524 3544 7530 3596
rect 7558 3544 7564 3596
rect 7616 3584 7622 3596
rect 8220 3593 8248 3624
rect 8294 3612 8300 3664
rect 8352 3652 8358 3664
rect 8352 3624 9260 3652
rect 8352 3612 8358 3624
rect 7929 3587 7987 3593
rect 7929 3584 7941 3587
rect 7616 3556 7941 3584
rect 7616 3544 7622 3556
rect 7929 3553 7941 3556
rect 7975 3553 7987 3587
rect 7929 3547 7987 3553
rect 8205 3587 8263 3593
rect 8205 3553 8217 3587
rect 8251 3553 8263 3587
rect 8386 3584 8392 3596
rect 8347 3556 8392 3584
rect 8205 3547 8263 3553
rect 8386 3544 8392 3556
rect 8444 3544 8450 3596
rect 8570 3584 8576 3596
rect 8483 3556 8576 3584
rect 8570 3544 8576 3556
rect 8628 3584 8634 3596
rect 9125 3587 9183 3593
rect 9125 3584 9137 3587
rect 8628 3556 9137 3584
rect 8628 3544 8634 3556
rect 9125 3553 9137 3556
rect 9171 3553 9183 3587
rect 9232 3584 9260 3624
rect 9692 3593 9720 3692
rect 10134 3680 10140 3692
rect 10192 3720 10198 3732
rect 10505 3723 10563 3729
rect 10505 3720 10517 3723
rect 10192 3692 10517 3720
rect 10192 3680 10198 3692
rect 10505 3689 10517 3692
rect 10551 3689 10563 3723
rect 10505 3683 10563 3689
rect 11054 3680 11060 3732
rect 11112 3680 11118 3732
rect 12710 3720 12716 3732
rect 11440 3692 12716 3720
rect 11072 3652 11100 3680
rect 10152 3624 11100 3652
rect 10152 3593 10180 3624
rect 9309 3587 9367 3593
rect 9309 3584 9321 3587
rect 9232 3556 9321 3584
rect 9125 3547 9183 3553
rect 9309 3553 9321 3556
rect 9355 3553 9367 3587
rect 9309 3547 9367 3553
rect 9677 3587 9735 3593
rect 9677 3553 9689 3587
rect 9723 3553 9735 3587
rect 9677 3547 9735 3553
rect 9953 3587 10011 3593
rect 9953 3553 9965 3587
rect 9999 3553 10011 3587
rect 9953 3547 10011 3553
rect 10137 3587 10195 3593
rect 10137 3553 10149 3587
rect 10183 3553 10195 3587
rect 10594 3584 10600 3596
rect 10555 3556 10600 3584
rect 10137 3547 10195 3553
rect 5626 3516 5632 3528
rect 5184 3488 5632 3516
rect 4663 3485 4675 3488
rect 4617 3479 4675 3485
rect 5626 3476 5632 3488
rect 5684 3476 5690 3528
rect 7650 3516 7656 3528
rect 5736 3488 7656 3516
rect 5736 3448 5764 3488
rect 7650 3476 7656 3488
rect 7708 3476 7714 3528
rect 7745 3519 7803 3525
rect 7745 3485 7757 3519
rect 7791 3485 7803 3519
rect 7745 3479 7803 3485
rect 7837 3519 7895 3525
rect 7837 3485 7849 3519
rect 7883 3516 7895 3519
rect 8754 3516 8760 3528
rect 7883 3488 8760 3516
rect 7883 3485 7895 3488
rect 7837 3479 7895 3485
rect 4080 3420 5764 3448
rect 3973 3411 4031 3417
rect 5810 3408 5816 3460
rect 5868 3448 5874 3460
rect 7760 3448 7788 3479
rect 8754 3476 8760 3488
rect 8812 3476 8818 3528
rect 9217 3519 9275 3525
rect 9217 3485 9229 3519
rect 9263 3516 9275 3519
rect 9490 3516 9496 3528
rect 9263 3488 9496 3516
rect 9263 3485 9275 3488
rect 9217 3479 9275 3485
rect 9490 3476 9496 3488
rect 9548 3476 9554 3528
rect 8386 3448 8392 3460
rect 5868 3420 6500 3448
rect 7760 3420 8392 3448
rect 5868 3408 5874 3420
rect 5442 3340 5448 3392
rect 5500 3380 5506 3392
rect 6472 3389 6500 3420
rect 8386 3408 8392 3420
rect 8444 3408 8450 3460
rect 6089 3383 6147 3389
rect 6089 3380 6101 3383
rect 5500 3352 6101 3380
rect 5500 3340 5506 3352
rect 6089 3349 6101 3352
rect 6135 3349 6147 3383
rect 6089 3343 6147 3349
rect 6457 3383 6515 3389
rect 6457 3349 6469 3383
rect 6503 3380 6515 3383
rect 8938 3380 8944 3392
rect 6503 3352 8944 3380
rect 6503 3349 6515 3352
rect 6457 3343 6515 3349
rect 8938 3340 8944 3352
rect 8996 3340 9002 3392
rect 9306 3340 9312 3392
rect 9364 3380 9370 3392
rect 9968 3380 9996 3547
rect 10594 3544 10600 3556
rect 10652 3544 10658 3596
rect 10686 3544 10692 3596
rect 10744 3584 10750 3596
rect 10781 3587 10839 3593
rect 10781 3584 10793 3587
rect 10744 3556 10793 3584
rect 10744 3544 10750 3556
rect 10781 3553 10793 3556
rect 10827 3553 10839 3587
rect 10781 3547 10839 3553
rect 10962 3544 10968 3596
rect 11020 3584 11026 3596
rect 11146 3584 11152 3596
rect 11020 3556 11065 3584
rect 11107 3556 11152 3584
rect 11020 3544 11026 3556
rect 11146 3544 11152 3556
rect 11204 3544 11210 3596
rect 10873 3519 10931 3525
rect 10873 3485 10885 3519
rect 10919 3516 10931 3519
rect 11440 3516 11468 3692
rect 12710 3680 12716 3692
rect 12768 3680 12774 3732
rect 12802 3612 12808 3664
rect 12860 3612 12866 3664
rect 10919 3488 11468 3516
rect 10919 3485 10931 3488
rect 10873 3479 10931 3485
rect 11514 3476 11520 3528
rect 11572 3516 11578 3528
rect 11790 3516 11796 3528
rect 11572 3488 11617 3516
rect 11751 3488 11796 3516
rect 11572 3476 11578 3488
rect 11790 3476 11796 3488
rect 11848 3476 11854 3528
rect 12158 3476 12164 3528
rect 12216 3516 12222 3528
rect 13265 3519 13323 3525
rect 13265 3516 13277 3519
rect 12216 3488 13277 3516
rect 12216 3476 12222 3488
rect 13265 3485 13277 3488
rect 13311 3485 13323 3519
rect 13265 3479 13323 3485
rect 12894 3380 12900 3392
rect 9364 3352 12900 3380
rect 9364 3340 9370 3352
rect 12894 3340 12900 3352
rect 12952 3340 12958 3392
rect 1104 3290 13892 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 12246 3290
rect 12298 3238 12310 3290
rect 12362 3238 12374 3290
rect 12426 3238 12438 3290
rect 12490 3238 13892 3290
rect 1104 3216 13892 3238
rect 4433 3179 4491 3185
rect 4433 3145 4445 3179
rect 4479 3176 4491 3179
rect 4614 3176 4620 3188
rect 4479 3148 4620 3176
rect 4479 3145 4491 3148
rect 4433 3139 4491 3145
rect 4614 3136 4620 3148
rect 4672 3136 4678 3188
rect 5169 3179 5227 3185
rect 5169 3145 5181 3179
rect 5215 3176 5227 3179
rect 6546 3176 6552 3188
rect 5215 3148 6552 3176
rect 5215 3145 5227 3148
rect 5169 3139 5227 3145
rect 6546 3136 6552 3148
rect 6604 3136 6610 3188
rect 7193 3179 7251 3185
rect 7193 3145 7205 3179
rect 7239 3176 7251 3179
rect 7466 3176 7472 3188
rect 7239 3148 7472 3176
rect 7239 3145 7251 3148
rect 7193 3139 7251 3145
rect 7466 3136 7472 3148
rect 7524 3136 7530 3188
rect 7558 3136 7564 3188
rect 7616 3176 7622 3188
rect 7837 3179 7895 3185
rect 7837 3176 7849 3179
rect 7616 3148 7849 3176
rect 7616 3136 7622 3148
rect 7837 3145 7849 3148
rect 7883 3145 7895 3179
rect 7837 3139 7895 3145
rect 8386 3136 8392 3188
rect 8444 3176 8450 3188
rect 8444 3148 9812 3176
rect 8444 3136 8450 3148
rect 1946 3108 1952 3120
rect 1907 3080 1952 3108
rect 1946 3068 1952 3080
rect 2004 3068 2010 3120
rect 4985 3111 5043 3117
rect 4985 3077 4997 3111
rect 5031 3077 5043 3111
rect 5534 3108 5540 3120
rect 5495 3080 5540 3108
rect 4985 3071 5043 3077
rect 1578 3000 1584 3052
rect 1636 3040 1642 3052
rect 4062 3040 4068 3052
rect 1636 3012 1992 3040
rect 4023 3012 4068 3040
rect 1636 3000 1642 3012
rect 1394 2932 1400 2984
rect 1452 2972 1458 2984
rect 1670 2972 1676 2984
rect 1452 2944 1676 2972
rect 1452 2932 1458 2944
rect 1670 2932 1676 2944
rect 1728 2972 1734 2984
rect 1765 2975 1823 2981
rect 1765 2972 1777 2975
rect 1728 2944 1777 2972
rect 1728 2932 1734 2944
rect 1765 2941 1777 2944
rect 1811 2941 1823 2975
rect 1765 2935 1823 2941
rect 1964 2916 1992 3012
rect 4062 3000 4068 3012
rect 4120 3000 4126 3052
rect 5000 3040 5028 3071
rect 5534 3068 5540 3080
rect 5592 3068 5598 3120
rect 5626 3068 5632 3120
rect 5684 3108 5690 3120
rect 9306 3108 9312 3120
rect 5684 3080 8432 3108
rect 9267 3080 9312 3108
rect 5684 3068 5690 3080
rect 6641 3043 6699 3049
rect 6641 3040 6653 3043
rect 5000 3012 6653 3040
rect 6641 3009 6653 3012
rect 6687 3040 6699 3043
rect 6687 3012 7604 3040
rect 6687 3009 6699 3012
rect 6641 3003 6699 3009
rect 4341 2975 4399 2981
rect 4341 2972 4353 2975
rect 4080 2944 4353 2972
rect 1486 2864 1492 2916
rect 1544 2904 1550 2916
rect 1581 2907 1639 2913
rect 1581 2904 1593 2907
rect 1544 2876 1593 2904
rect 1544 2864 1550 2876
rect 1581 2873 1593 2876
rect 1627 2873 1639 2907
rect 1581 2867 1639 2873
rect 1946 2864 1952 2916
rect 2004 2904 2010 2916
rect 3786 2904 3792 2916
rect 2004 2876 2622 2904
rect 3747 2876 3792 2904
rect 2004 2864 2010 2876
rect 3786 2864 3792 2876
rect 3844 2864 3850 2916
rect 2317 2839 2375 2845
rect 2317 2805 2329 2839
rect 2363 2836 2375 2839
rect 2498 2836 2504 2848
rect 2363 2808 2504 2836
rect 2363 2805 2375 2808
rect 2317 2799 2375 2805
rect 2498 2796 2504 2808
rect 2556 2796 2562 2848
rect 3418 2796 3424 2848
rect 3476 2836 3482 2848
rect 4080 2836 4108 2944
rect 4341 2941 4353 2944
rect 4387 2941 4399 2975
rect 4341 2935 4399 2941
rect 4706 2932 4712 2984
rect 4764 2972 4770 2984
rect 4803 2975 4861 2981
rect 4803 2972 4815 2975
rect 4764 2944 4815 2972
rect 4764 2932 4770 2944
rect 4803 2941 4815 2944
rect 4849 2941 4861 2975
rect 4803 2935 4861 2941
rect 5169 2975 5227 2981
rect 5169 2941 5181 2975
rect 5215 2972 5227 2975
rect 5353 2975 5411 2981
rect 5353 2972 5365 2975
rect 5215 2944 5365 2972
rect 5215 2941 5227 2944
rect 5169 2935 5227 2941
rect 5353 2941 5365 2944
rect 5399 2941 5411 2975
rect 5353 2935 5411 2941
rect 5721 2975 5779 2981
rect 5721 2941 5733 2975
rect 5767 2941 5779 2975
rect 5902 2972 5908 2984
rect 5863 2944 5908 2972
rect 5721 2935 5779 2941
rect 4798 2836 4804 2848
rect 3476 2808 4108 2836
rect 4759 2808 4804 2836
rect 3476 2796 3482 2808
rect 4798 2796 4804 2808
rect 4856 2796 4862 2848
rect 5736 2836 5764 2935
rect 5902 2932 5908 2944
rect 5960 2972 5966 2984
rect 6270 2972 6276 2984
rect 5960 2944 6276 2972
rect 5960 2932 5966 2944
rect 6270 2932 6276 2944
rect 6328 2932 6334 2984
rect 6730 2972 6736 2984
rect 6691 2944 6736 2972
rect 6730 2932 6736 2944
rect 6788 2932 6794 2984
rect 7576 2981 7604 3012
rect 7071 2975 7129 2981
rect 7071 2941 7083 2975
rect 7117 2972 7129 2975
rect 7469 2975 7527 2981
rect 7469 2972 7481 2975
rect 7117 2944 7481 2972
rect 7117 2941 7129 2944
rect 7071 2935 7129 2941
rect 7469 2941 7481 2944
rect 7515 2941 7527 2975
rect 7469 2935 7527 2941
rect 7561 2975 7619 2981
rect 7561 2941 7573 2975
rect 7607 2941 7619 2975
rect 7561 2935 7619 2941
rect 7650 2932 7656 2984
rect 7708 2972 7714 2984
rect 8404 2981 8432 3080
rect 9306 3068 9312 3080
rect 9364 3068 9370 3120
rect 9784 3108 9812 3148
rect 9858 3136 9864 3188
rect 9916 3176 9922 3188
rect 10781 3179 10839 3185
rect 10781 3176 10793 3179
rect 9916 3148 10793 3176
rect 9916 3136 9922 3148
rect 10781 3145 10793 3148
rect 10827 3145 10839 3179
rect 10781 3139 10839 3145
rect 11054 3136 11060 3188
rect 11112 3176 11118 3188
rect 11425 3179 11483 3185
rect 11425 3176 11437 3179
rect 11112 3148 11437 3176
rect 11112 3136 11118 3148
rect 11425 3145 11437 3148
rect 11471 3145 11483 3179
rect 11790 3176 11796 3188
rect 11751 3148 11796 3176
rect 11425 3139 11483 3145
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 12621 3179 12679 3185
rect 12621 3145 12633 3179
rect 12667 3176 12679 3179
rect 12802 3176 12808 3188
rect 12667 3148 12808 3176
rect 12667 3145 12679 3148
rect 12621 3139 12679 3145
rect 12802 3136 12808 3148
rect 12860 3136 12866 3188
rect 12986 3136 12992 3188
rect 13044 3176 13050 3188
rect 13081 3179 13139 3185
rect 13081 3176 13093 3179
rect 13044 3148 13093 3176
rect 13044 3136 13050 3148
rect 13081 3145 13093 3148
rect 13127 3145 13139 3179
rect 13081 3139 13139 3145
rect 12526 3108 12532 3120
rect 9784 3080 12532 3108
rect 12526 3068 12532 3080
rect 12584 3068 12590 3120
rect 9398 3040 9404 3052
rect 9311 3012 9404 3040
rect 9398 3000 9404 3012
rect 9456 3040 9462 3052
rect 11238 3040 11244 3052
rect 9456 3012 10180 3040
rect 9456 3000 9462 3012
rect 8205 2975 8263 2981
rect 8205 2972 8217 2975
rect 7708 2944 8217 2972
rect 7708 2932 7714 2944
rect 8205 2941 8217 2944
rect 8251 2941 8263 2975
rect 8205 2935 8263 2941
rect 8389 2975 8447 2981
rect 8389 2941 8401 2975
rect 8435 2941 8447 2975
rect 8846 2972 8852 2984
rect 8807 2944 8852 2972
rect 8389 2935 8447 2941
rect 8846 2932 8852 2944
rect 8904 2932 8910 2984
rect 8938 2932 8944 2984
rect 8996 2972 9002 2984
rect 9033 2975 9091 2981
rect 9033 2972 9045 2975
rect 8996 2944 9045 2972
rect 8996 2932 9002 2944
rect 9033 2941 9045 2944
rect 9079 2941 9091 2975
rect 9033 2935 9091 2941
rect 9122 2932 9128 2984
rect 9180 2972 9186 2984
rect 9950 2981 9956 2984
rect 9752 2975 9810 2981
rect 9752 2972 9764 2975
rect 9180 2944 9764 2972
rect 9180 2932 9186 2944
rect 9752 2941 9764 2944
rect 9798 2941 9810 2975
rect 9752 2935 9810 2941
rect 9948 2935 9956 2981
rect 10008 2972 10014 2984
rect 10152 2981 10180 3012
rect 11072 3012 11244 3040
rect 10137 2975 10195 2981
rect 10008 2944 10048 2972
rect 9950 2932 9956 2935
rect 10008 2932 10014 2944
rect 10137 2941 10149 2975
rect 10183 2941 10195 2975
rect 10318 2972 10324 2984
rect 10279 2944 10324 2972
rect 10137 2935 10195 2941
rect 10318 2932 10324 2944
rect 10376 2932 10382 2984
rect 11072 2981 11100 3012
rect 11238 3000 11244 3012
rect 11296 3000 11302 3052
rect 11698 3000 11704 3052
rect 11756 3040 11762 3052
rect 11756 3012 12388 3040
rect 11756 3000 11762 3012
rect 11057 2975 11115 2981
rect 11057 2941 11069 2975
rect 11103 2941 11115 2975
rect 11057 2935 11115 2941
rect 11149 2975 11207 2981
rect 11149 2941 11161 2975
rect 11195 2972 11207 2975
rect 11425 2975 11483 2981
rect 11425 2972 11437 2975
rect 11195 2944 11437 2972
rect 11195 2941 11207 2944
rect 11149 2935 11207 2941
rect 11425 2941 11437 2944
rect 11471 2972 11483 2975
rect 11716 2972 11744 3000
rect 11471 2944 11744 2972
rect 11471 2941 11483 2944
rect 11425 2935 11483 2941
rect 11882 2932 11888 2984
rect 11940 2981 11946 2984
rect 12360 2981 12388 3012
rect 11940 2975 11983 2981
rect 11971 2941 11983 2975
rect 11940 2935 11983 2941
rect 12345 2975 12403 2981
rect 12345 2941 12357 2975
rect 12391 2941 12403 2975
rect 12802 2972 12808 2984
rect 12763 2944 12808 2972
rect 12345 2935 12403 2941
rect 11940 2932 11946 2935
rect 12802 2932 12808 2944
rect 12860 2972 12866 2984
rect 13078 2972 13084 2984
rect 12860 2944 13084 2972
rect 12860 2932 12866 2944
rect 13078 2932 13084 2944
rect 13136 2932 13142 2984
rect 13262 2972 13268 2984
rect 13223 2944 13268 2972
rect 13262 2932 13268 2944
rect 13320 2932 13326 2984
rect 6748 2904 6776 2932
rect 7745 2907 7803 2913
rect 7745 2904 7757 2907
rect 6748 2876 7757 2904
rect 7745 2873 7757 2876
rect 7791 2873 7803 2907
rect 8570 2904 8576 2916
rect 8531 2876 8576 2904
rect 7745 2867 7803 2873
rect 8570 2864 8576 2876
rect 8628 2864 8634 2916
rect 10045 2907 10103 2913
rect 10045 2873 10057 2907
rect 10091 2873 10103 2907
rect 10045 2867 10103 2873
rect 11333 2907 11391 2913
rect 11333 2873 11345 2907
rect 11379 2904 11391 2907
rect 12066 2904 12072 2916
rect 11379 2876 12072 2904
rect 11379 2873 11391 2876
rect 11333 2867 11391 2873
rect 5810 2836 5816 2848
rect 5736 2808 5816 2836
rect 5810 2796 5816 2808
rect 5868 2796 5874 2848
rect 10060 2836 10088 2867
rect 12066 2864 12072 2876
rect 12124 2864 12130 2916
rect 12161 2907 12219 2913
rect 12161 2873 12173 2907
rect 12207 2873 12219 2907
rect 12161 2867 12219 2873
rect 10226 2836 10232 2848
rect 10060 2808 10232 2836
rect 10226 2796 10232 2808
rect 10284 2796 10290 2848
rect 10965 2839 11023 2845
rect 10965 2805 10977 2839
rect 11011 2836 11023 2839
rect 11238 2836 11244 2848
rect 11011 2808 11244 2836
rect 11011 2805 11023 2808
rect 10965 2799 11023 2805
rect 11238 2796 11244 2808
rect 11296 2836 11302 2848
rect 12176 2836 12204 2867
rect 12250 2836 12256 2848
rect 11296 2808 12256 2836
rect 11296 2796 11302 2808
rect 12250 2796 12256 2808
rect 12308 2796 12314 2848
rect 1104 2746 13892 2768
rect 1104 2694 8246 2746
rect 8298 2694 8310 2746
rect 8362 2694 8374 2746
rect 8426 2694 8438 2746
rect 8490 2694 13892 2746
rect 1104 2672 13892 2694
rect 2041 2635 2099 2641
rect 2041 2601 2053 2635
rect 2087 2632 2099 2635
rect 4614 2632 4620 2644
rect 2087 2604 4620 2632
rect 2087 2601 2099 2604
rect 2041 2595 2099 2601
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 5350 2632 5356 2644
rect 5311 2604 5356 2632
rect 5350 2592 5356 2604
rect 5408 2592 5414 2644
rect 5537 2635 5595 2641
rect 5537 2601 5549 2635
rect 5583 2632 5595 2635
rect 5626 2632 5632 2644
rect 5583 2604 5632 2632
rect 5583 2601 5595 2604
rect 5537 2595 5595 2601
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 6362 2632 6368 2644
rect 5736 2604 6368 2632
rect 3050 2564 3056 2576
rect 3011 2536 3056 2564
rect 3050 2524 3056 2536
rect 3108 2524 3114 2576
rect 3513 2567 3571 2573
rect 3513 2564 3525 2567
rect 3160 2536 3525 2564
rect 1857 2499 1915 2505
rect 1857 2465 1869 2499
rect 1903 2496 1915 2499
rect 1946 2496 1952 2508
rect 1903 2468 1952 2496
rect 1903 2465 1915 2468
rect 1857 2459 1915 2465
rect 1946 2456 1952 2468
rect 2004 2456 2010 2508
rect 2314 2496 2320 2508
rect 2275 2468 2320 2496
rect 2314 2456 2320 2468
rect 2372 2456 2378 2508
rect 2498 2496 2504 2508
rect 2459 2468 2504 2496
rect 2498 2456 2504 2468
rect 2556 2496 2562 2508
rect 3160 2496 3188 2536
rect 3513 2533 3525 2536
rect 3559 2564 3571 2567
rect 4249 2567 4307 2573
rect 4249 2564 4261 2567
rect 3559 2536 4261 2564
rect 3559 2533 3571 2536
rect 3513 2527 3571 2533
rect 4249 2533 4261 2536
rect 4295 2564 4307 2567
rect 4798 2564 4804 2576
rect 4295 2536 4804 2564
rect 4295 2533 4307 2536
rect 4249 2527 4307 2533
rect 4798 2524 4804 2536
rect 4856 2524 4862 2576
rect 5261 2567 5319 2573
rect 5261 2533 5273 2567
rect 5307 2564 5319 2567
rect 5736 2564 5764 2604
rect 6362 2592 6368 2604
rect 6420 2592 6426 2644
rect 7101 2635 7159 2641
rect 7101 2601 7113 2635
rect 7147 2632 7159 2635
rect 7650 2632 7656 2644
rect 7147 2604 7656 2632
rect 7147 2601 7159 2604
rect 7101 2595 7159 2601
rect 7650 2592 7656 2604
rect 7708 2592 7714 2644
rect 10505 2635 10563 2641
rect 10505 2632 10517 2635
rect 8128 2604 10517 2632
rect 5307 2536 5764 2564
rect 5307 2533 5319 2536
rect 5261 2527 5319 2533
rect 5644 2508 5672 2536
rect 6270 2524 6276 2576
rect 6328 2564 6334 2576
rect 7929 2567 7987 2573
rect 7929 2564 7941 2567
rect 6328 2536 7052 2564
rect 6328 2524 6334 2536
rect 2556 2468 3188 2496
rect 3237 2499 3295 2505
rect 2556 2456 2562 2468
rect 3237 2465 3249 2499
rect 3283 2496 3295 2499
rect 3326 2496 3332 2508
rect 3283 2468 3332 2496
rect 3283 2465 3295 2468
rect 3237 2459 3295 2465
rect 2685 2431 2743 2437
rect 2685 2397 2697 2431
rect 2731 2428 2743 2431
rect 3252 2428 3280 2459
rect 3326 2456 3332 2468
rect 3384 2456 3390 2508
rect 4154 2505 4160 2508
rect 3421 2499 3479 2505
rect 3421 2465 3433 2499
rect 3467 2465 3479 2499
rect 4152 2496 4160 2505
rect 4115 2468 4160 2496
rect 3421 2459 3479 2465
rect 4152 2459 4160 2468
rect 2731 2400 3280 2428
rect 3436 2428 3464 2459
rect 4154 2456 4160 2459
rect 4212 2456 4218 2508
rect 4341 2499 4399 2505
rect 4341 2465 4353 2499
rect 4387 2465 4399 2499
rect 4341 2459 4399 2465
rect 4525 2499 4583 2505
rect 4525 2465 4537 2499
rect 4571 2496 4583 2499
rect 5166 2496 5172 2508
rect 4571 2468 5028 2496
rect 5127 2468 5172 2496
rect 4571 2465 4583 2468
rect 4525 2459 4583 2465
rect 4356 2428 4384 2459
rect 5000 2428 5028 2468
rect 5166 2456 5172 2468
rect 5224 2456 5230 2508
rect 5350 2456 5356 2508
rect 5408 2496 5414 2508
rect 5408 2468 5580 2496
rect 5408 2456 5414 2468
rect 5552 2428 5580 2468
rect 5626 2456 5632 2508
rect 5684 2456 5690 2508
rect 6178 2496 6184 2508
rect 6139 2468 6184 2496
rect 6178 2456 6184 2468
rect 6236 2456 6242 2508
rect 6457 2499 6515 2505
rect 6457 2465 6469 2499
rect 6503 2465 6515 2499
rect 6457 2459 6515 2465
rect 6365 2431 6423 2437
rect 6365 2428 6377 2431
rect 3436 2400 4660 2428
rect 5000 2400 5304 2428
rect 5552 2400 6377 2428
rect 2731 2397 2743 2400
rect 2685 2391 2743 2397
rect 2314 2320 2320 2372
rect 2372 2360 2378 2372
rect 3326 2360 3332 2372
rect 2372 2332 3332 2360
rect 2372 2320 2378 2332
rect 3326 2320 3332 2332
rect 3384 2360 3390 2372
rect 3436 2360 3464 2400
rect 4632 2372 4660 2400
rect 3384 2332 3464 2360
rect 3384 2320 3390 2332
rect 3786 2320 3792 2372
rect 3844 2360 3850 2372
rect 3973 2363 4031 2369
rect 3973 2360 3985 2363
rect 3844 2332 3985 2360
rect 3844 2320 3850 2332
rect 3973 2329 3985 2332
rect 4019 2329 4031 2363
rect 3973 2323 4031 2329
rect 4154 2320 4160 2372
rect 4212 2320 4218 2372
rect 4614 2320 4620 2372
rect 4672 2360 4678 2372
rect 4985 2363 5043 2369
rect 4985 2360 4997 2363
rect 4672 2332 4997 2360
rect 4672 2320 4678 2332
rect 4985 2329 4997 2332
rect 5031 2329 5043 2363
rect 5276 2360 5304 2400
rect 6365 2397 6377 2400
rect 6411 2428 6423 2431
rect 6472 2428 6500 2459
rect 6546 2456 6552 2508
rect 6604 2505 6610 2508
rect 6604 2499 6663 2505
rect 6604 2465 6617 2499
rect 6651 2465 6663 2499
rect 6604 2459 6663 2465
rect 6604 2456 6610 2459
rect 6730 2456 6736 2508
rect 6788 2496 6794 2508
rect 7024 2505 7052 2536
rect 7116 2536 7941 2564
rect 7009 2499 7067 2505
rect 6788 2468 6960 2496
rect 6788 2456 6794 2468
rect 6411 2400 6500 2428
rect 6825 2431 6883 2437
rect 6411 2397 6423 2400
rect 6365 2391 6423 2397
rect 6825 2397 6837 2431
rect 6871 2397 6883 2431
rect 6932 2428 6960 2468
rect 7009 2465 7021 2499
rect 7055 2465 7067 2499
rect 7009 2459 7067 2465
rect 7116 2428 7144 2536
rect 7929 2533 7941 2536
rect 7975 2533 7987 2567
rect 7929 2527 7987 2533
rect 8128 2508 8156 2604
rect 10505 2601 10517 2604
rect 10551 2601 10563 2635
rect 10686 2632 10692 2644
rect 10505 2595 10563 2601
rect 10612 2604 10692 2632
rect 8938 2564 8944 2576
rect 8496 2536 8944 2564
rect 7740 2499 7798 2505
rect 7740 2465 7752 2499
rect 7786 2465 7798 2499
rect 7740 2459 7798 2465
rect 7837 2499 7895 2505
rect 7837 2465 7849 2499
rect 7883 2465 7895 2499
rect 8110 2496 8116 2508
rect 8071 2468 8116 2496
rect 7837 2459 7895 2465
rect 6932 2400 7144 2428
rect 6825 2391 6883 2397
rect 5718 2360 5724 2372
rect 5276 2332 5724 2360
rect 4985 2323 5043 2329
rect 5718 2320 5724 2332
rect 5776 2320 5782 2372
rect 5810 2320 5816 2372
rect 5868 2360 5874 2372
rect 6638 2360 6644 2372
rect 5868 2332 6644 2360
rect 5868 2320 5874 2332
rect 6638 2320 6644 2332
rect 6696 2360 6702 2372
rect 6840 2360 6868 2391
rect 7760 2360 7788 2459
rect 7852 2428 7880 2459
rect 8110 2456 8116 2468
rect 8168 2456 8174 2508
rect 8496 2505 8524 2536
rect 8938 2524 8944 2536
rect 8996 2524 9002 2576
rect 9861 2567 9919 2573
rect 9861 2533 9873 2567
rect 9907 2564 9919 2567
rect 10612 2564 10640 2604
rect 10686 2592 10692 2604
rect 10744 2592 10750 2644
rect 12250 2592 12256 2644
rect 12308 2632 12314 2644
rect 13081 2635 13139 2641
rect 13081 2632 13093 2635
rect 12308 2604 13093 2632
rect 12308 2592 12314 2604
rect 13081 2601 13093 2604
rect 13127 2601 13139 2635
rect 13081 2595 13139 2601
rect 9907 2536 10640 2564
rect 9907 2533 9919 2536
rect 9861 2527 9919 2533
rect 8481 2499 8539 2505
rect 8481 2465 8493 2499
rect 8527 2465 8539 2499
rect 8481 2459 8539 2465
rect 8665 2499 8723 2505
rect 8665 2465 8677 2499
rect 8711 2496 8723 2499
rect 8846 2496 8852 2508
rect 8711 2468 8852 2496
rect 8711 2465 8723 2468
rect 8665 2459 8723 2465
rect 8846 2456 8852 2468
rect 8904 2496 8910 2508
rect 9214 2496 9220 2508
rect 8904 2468 9220 2496
rect 8904 2456 8910 2468
rect 9214 2456 9220 2468
rect 9272 2456 9278 2508
rect 9493 2499 9551 2505
rect 9493 2465 9505 2499
rect 9539 2496 9551 2499
rect 10137 2499 10195 2505
rect 10137 2496 10149 2499
rect 9539 2468 10149 2496
rect 9539 2465 9551 2468
rect 9493 2459 9551 2465
rect 10137 2465 10149 2468
rect 10183 2496 10195 2499
rect 10318 2496 10324 2508
rect 10183 2468 10324 2496
rect 10183 2465 10195 2468
rect 10137 2459 10195 2465
rect 10318 2456 10324 2468
rect 10376 2456 10382 2508
rect 10612 2505 10640 2536
rect 10965 2567 11023 2573
rect 10965 2533 10977 2567
rect 11011 2564 11023 2567
rect 11146 2564 11152 2576
rect 11011 2536 11152 2564
rect 11011 2533 11023 2536
rect 10965 2527 11023 2533
rect 11146 2524 11152 2536
rect 11204 2524 11210 2576
rect 11514 2564 11520 2576
rect 11348 2536 11520 2564
rect 10597 2499 10655 2505
rect 10597 2465 10609 2499
rect 10643 2465 10655 2499
rect 10597 2459 10655 2465
rect 10686 2456 10692 2508
rect 10744 2496 10750 2508
rect 11348 2505 11376 2536
rect 11514 2524 11520 2536
rect 11572 2524 11578 2576
rect 12618 2524 12624 2576
rect 12676 2524 12682 2576
rect 10781 2499 10839 2505
rect 10781 2496 10793 2499
rect 10744 2468 10793 2496
rect 10744 2456 10750 2468
rect 10781 2465 10793 2468
rect 10827 2465 10839 2499
rect 10781 2459 10839 2465
rect 11333 2499 11391 2505
rect 11333 2465 11345 2499
rect 11379 2465 11391 2499
rect 11333 2459 11391 2465
rect 8754 2428 8760 2440
rect 7852 2400 8760 2428
rect 8754 2388 8760 2400
rect 8812 2388 8818 2440
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2428 9367 2431
rect 9398 2428 9404 2440
rect 9355 2400 9404 2428
rect 9355 2397 9367 2400
rect 9309 2391 9367 2397
rect 8665 2363 8723 2369
rect 6696 2332 6868 2360
rect 7392 2332 8294 2360
rect 6696 2320 6702 2332
rect 4172 2292 4200 2320
rect 5350 2292 5356 2304
rect 4172 2264 5356 2292
rect 5350 2252 5356 2264
rect 5408 2252 5414 2304
rect 5534 2252 5540 2304
rect 5592 2292 5598 2304
rect 5997 2295 6055 2301
rect 5997 2292 6009 2295
rect 5592 2264 6009 2292
rect 5592 2252 5598 2264
rect 5997 2261 6009 2264
rect 6043 2261 6055 2295
rect 5997 2255 6055 2261
rect 6365 2295 6423 2301
rect 6365 2261 6377 2295
rect 6411 2292 6423 2295
rect 7392 2292 7420 2332
rect 7558 2292 7564 2304
rect 6411 2264 7420 2292
rect 7519 2264 7564 2292
rect 6411 2261 6423 2264
rect 6365 2255 6423 2261
rect 7558 2252 7564 2264
rect 7616 2252 7622 2304
rect 8266 2292 8294 2332
rect 8665 2329 8677 2363
rect 8711 2360 8723 2363
rect 9324 2360 9352 2391
rect 9398 2388 9404 2400
rect 9456 2428 9462 2440
rect 10045 2431 10103 2437
rect 10045 2428 10057 2431
rect 9456 2400 10057 2428
rect 9456 2388 9462 2400
rect 10045 2397 10057 2400
rect 10091 2397 10103 2431
rect 11606 2428 11612 2440
rect 11567 2400 11612 2428
rect 10045 2391 10103 2397
rect 11606 2388 11612 2400
rect 11664 2388 11670 2440
rect 8711 2332 9352 2360
rect 10505 2363 10563 2369
rect 8711 2329 8723 2332
rect 8665 2323 8723 2329
rect 10505 2329 10517 2363
rect 10551 2360 10563 2363
rect 11054 2360 11060 2372
rect 10551 2332 11060 2360
rect 10551 2329 10563 2332
rect 10505 2323 10563 2329
rect 11054 2320 11060 2332
rect 11112 2320 11118 2372
rect 11790 2292 11796 2304
rect 8266 2264 11796 2292
rect 11790 2252 11796 2264
rect 11848 2252 11854 2304
rect 1104 2202 13892 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 12246 2202
rect 12298 2150 12310 2202
rect 12362 2150 12374 2202
rect 12426 2150 12438 2202
rect 12490 2150 13892 2202
rect 1104 2128 13892 2150
rect 2133 2091 2191 2097
rect 2133 2057 2145 2091
rect 2179 2088 2191 2091
rect 2314 2088 2320 2100
rect 2179 2060 2320 2088
rect 2179 2057 2191 2060
rect 2133 2051 2191 2057
rect 2314 2048 2320 2060
rect 2372 2048 2378 2100
rect 4614 2048 4620 2100
rect 4672 2088 4678 2100
rect 4672 2060 5764 2088
rect 4672 2048 4678 2060
rect 4246 1980 4252 2032
rect 4304 2020 4310 2032
rect 5442 2020 5448 2032
rect 4304 1992 5448 2020
rect 4304 1980 4310 1992
rect 5442 1980 5448 1992
rect 5500 1980 5506 2032
rect 3881 1955 3939 1961
rect 3881 1921 3893 1955
rect 3927 1952 3939 1955
rect 4062 1952 4068 1964
rect 3927 1924 4068 1952
rect 3927 1921 3939 1924
rect 3881 1915 3939 1921
rect 4062 1912 4068 1924
rect 4120 1912 4126 1964
rect 4154 1912 4160 1964
rect 4212 1952 4218 1964
rect 4798 1952 4804 1964
rect 4212 1924 4804 1952
rect 4212 1912 4218 1924
rect 4798 1912 4804 1924
rect 4856 1912 4862 1964
rect 4908 1924 5672 1952
rect 4525 1887 4583 1893
rect 4525 1853 4537 1887
rect 4571 1884 4583 1887
rect 4614 1884 4620 1896
rect 4571 1856 4620 1884
rect 4571 1853 4583 1856
rect 4525 1847 4583 1853
rect 4614 1844 4620 1856
rect 4672 1844 4678 1896
rect 4908 1893 4936 1924
rect 5644 1896 5672 1924
rect 4709 1887 4767 1893
rect 4709 1853 4721 1887
rect 4755 1853 4767 1887
rect 4709 1847 4767 1853
rect 4894 1887 4952 1893
rect 4894 1853 4906 1887
rect 4940 1853 4952 1887
rect 4894 1847 4952 1853
rect 5077 1887 5135 1893
rect 5077 1853 5089 1887
rect 5123 1884 5135 1887
rect 5350 1884 5356 1896
rect 5123 1856 5356 1884
rect 5123 1853 5135 1856
rect 5077 1847 5135 1853
rect 2866 1776 2872 1828
rect 2924 1776 2930 1828
rect 3605 1819 3663 1825
rect 3605 1785 3617 1819
rect 3651 1816 3663 1819
rect 4341 1819 4399 1825
rect 4341 1816 4353 1819
rect 3651 1788 4353 1816
rect 3651 1785 3663 1788
rect 3605 1779 3663 1785
rect 4341 1785 4353 1788
rect 4387 1785 4399 1819
rect 4724 1816 4752 1847
rect 5350 1844 5356 1856
rect 5408 1844 5414 1896
rect 5626 1884 5632 1896
rect 5587 1856 5632 1884
rect 5626 1844 5632 1856
rect 5684 1844 5690 1896
rect 5736 1884 5764 2060
rect 6270 2048 6276 2100
rect 6328 2088 6334 2100
rect 6641 2091 6699 2097
rect 6641 2088 6653 2091
rect 6328 2060 6653 2088
rect 6328 2048 6334 2060
rect 6641 2057 6653 2060
rect 6687 2057 6699 2091
rect 6641 2051 6699 2057
rect 7101 2091 7159 2097
rect 7101 2057 7113 2091
rect 7147 2088 7159 2091
rect 9214 2088 9220 2100
rect 7147 2060 9076 2088
rect 9175 2060 9220 2088
rect 7147 2057 7159 2060
rect 7101 2051 7159 2057
rect 5810 1912 5816 1964
rect 5868 1952 5874 1964
rect 5868 1924 5948 1952
rect 5868 1912 5874 1924
rect 5920 1893 5948 1924
rect 5905 1887 5963 1893
rect 5736 1856 5856 1884
rect 5166 1816 5172 1828
rect 4341 1779 4399 1785
rect 4540 1788 5172 1816
rect 3970 1708 3976 1760
rect 4028 1748 4034 1760
rect 4540 1748 4568 1788
rect 5166 1776 5172 1788
rect 5224 1816 5230 1828
rect 5828 1825 5856 1856
rect 5905 1853 5917 1887
rect 5951 1853 5963 1887
rect 5905 1847 5963 1853
rect 5994 1844 6000 1896
rect 6052 1884 6058 1896
rect 6089 1887 6147 1893
rect 6089 1884 6101 1887
rect 6052 1856 6101 1884
rect 6052 1844 6058 1856
rect 6089 1853 6101 1856
rect 6135 1853 6147 1887
rect 6089 1847 6147 1853
rect 5721 1819 5779 1825
rect 5721 1816 5733 1819
rect 5224 1788 5733 1816
rect 5224 1776 5230 1788
rect 5721 1785 5733 1788
rect 5767 1785 5779 1819
rect 5721 1779 5779 1785
rect 5813 1819 5871 1825
rect 5813 1785 5825 1819
rect 5859 1785 5871 1819
rect 6104 1816 6132 1847
rect 6546 1844 6552 1896
rect 6604 1884 6610 1896
rect 6733 1887 6791 1893
rect 6733 1884 6745 1887
rect 6604 1856 6745 1884
rect 6604 1844 6610 1856
rect 6733 1853 6745 1856
rect 6779 1884 6791 1887
rect 7116 1884 7144 2051
rect 9048 2020 9076 2060
rect 9214 2048 9220 2060
rect 9272 2048 9278 2100
rect 9861 2091 9919 2097
rect 9861 2057 9873 2091
rect 9907 2088 9919 2091
rect 10318 2088 10324 2100
rect 9907 2060 10324 2088
rect 9907 2057 9919 2060
rect 9861 2051 9919 2057
rect 10318 2048 10324 2060
rect 10376 2048 10382 2100
rect 11241 2091 11299 2097
rect 11241 2057 11253 2091
rect 11287 2088 11299 2091
rect 11606 2088 11612 2100
rect 11287 2060 11612 2088
rect 11287 2057 11299 2060
rect 11241 2051 11299 2057
rect 11606 2048 11612 2060
rect 11664 2048 11670 2100
rect 12710 2048 12716 2100
rect 12768 2088 12774 2100
rect 13173 2091 13231 2097
rect 13173 2088 13185 2091
rect 12768 2060 13185 2088
rect 12768 2048 12774 2060
rect 13173 2057 13185 2060
rect 13219 2057 13231 2091
rect 13173 2051 13231 2057
rect 9048 1992 9260 2020
rect 8110 1952 8116 1964
rect 6779 1856 7144 1884
rect 7300 1924 8116 1952
rect 6779 1853 6791 1856
rect 6733 1847 6791 1853
rect 7300 1816 7328 1924
rect 8110 1912 8116 1924
rect 8168 1912 8174 1964
rect 8570 1952 8576 1964
rect 8531 1924 8576 1952
rect 8570 1912 8576 1924
rect 8628 1912 8634 1964
rect 8849 1955 8907 1961
rect 8849 1921 8861 1955
rect 8895 1952 8907 1955
rect 9033 1955 9091 1961
rect 9033 1952 9045 1955
rect 8895 1924 9045 1952
rect 8895 1921 8907 1924
rect 8849 1915 8907 1921
rect 9033 1921 9045 1924
rect 9079 1921 9091 1955
rect 9033 1915 9091 1921
rect 8938 1844 8944 1896
rect 8996 1884 9002 1896
rect 9125 1887 9183 1893
rect 9125 1884 9137 1887
rect 8996 1856 9137 1884
rect 8996 1844 9002 1856
rect 9125 1853 9137 1856
rect 9171 1853 9183 1887
rect 9232 1884 9260 1992
rect 10042 1980 10048 2032
rect 10100 2020 10106 2032
rect 10413 2023 10471 2029
rect 10413 2020 10425 2023
rect 10100 1992 10425 2020
rect 10100 1980 10106 1992
rect 10413 1989 10425 1992
rect 10459 1989 10471 2023
rect 10413 1983 10471 1989
rect 10428 1952 10456 1983
rect 11054 1980 11060 2032
rect 11112 2020 11118 2032
rect 11517 2023 11575 2029
rect 11517 2020 11529 2023
rect 11112 1992 11529 2020
rect 11112 1980 11118 1992
rect 11517 1989 11529 1992
rect 11563 1989 11575 2023
rect 11517 1983 11575 1989
rect 11882 1980 11888 2032
rect 11940 2020 11946 2032
rect 12250 2020 12256 2032
rect 11940 1992 12112 2020
rect 12211 1992 12256 2020
rect 11940 1980 11946 1992
rect 10428 1924 12020 1952
rect 10043 1887 10101 1893
rect 10043 1884 10055 1887
rect 9232 1856 10055 1884
rect 9125 1847 9183 1853
rect 10043 1853 10055 1856
rect 10089 1884 10101 1887
rect 10226 1884 10232 1896
rect 10089 1856 10232 1884
rect 10089 1853 10101 1856
rect 10043 1847 10101 1853
rect 10226 1844 10232 1856
rect 10284 1884 10290 1896
rect 10505 1887 10563 1893
rect 10505 1884 10517 1887
rect 10284 1856 10517 1884
rect 10284 1844 10290 1856
rect 10505 1853 10517 1856
rect 10551 1884 10563 1887
rect 11149 1887 11207 1893
rect 10551 1856 11100 1884
rect 10551 1853 10563 1856
rect 10505 1847 10563 1853
rect 10962 1816 10968 1828
rect 6104 1788 7328 1816
rect 8142 1788 10272 1816
rect 10923 1788 10968 1816
rect 5813 1779 5871 1785
rect 4028 1720 4568 1748
rect 4028 1708 4034 1720
rect 4614 1708 4620 1760
rect 4672 1748 4678 1760
rect 5445 1751 5503 1757
rect 5445 1748 5457 1751
rect 4672 1720 5457 1748
rect 4672 1708 4678 1720
rect 5445 1717 5457 1720
rect 5491 1717 5503 1751
rect 5445 1711 5503 1717
rect 6178 1708 6184 1760
rect 6236 1748 6242 1760
rect 6822 1748 6828 1760
rect 6236 1720 6828 1748
rect 6236 1708 6242 1720
rect 6822 1708 6828 1720
rect 6880 1748 6886 1760
rect 9033 1751 9091 1757
rect 9033 1748 9045 1751
rect 6880 1720 9045 1748
rect 6880 1708 6886 1720
rect 9033 1717 9045 1720
rect 9079 1717 9091 1751
rect 9033 1711 9091 1717
rect 9766 1708 9772 1760
rect 9824 1748 9830 1760
rect 10042 1748 10048 1760
rect 9824 1720 10048 1748
rect 9824 1708 9830 1720
rect 10042 1708 10048 1720
rect 10100 1708 10106 1760
rect 10244 1748 10272 1788
rect 10962 1776 10968 1788
rect 11020 1776 11026 1828
rect 11072 1816 11100 1856
rect 11149 1853 11161 1887
rect 11195 1884 11207 1887
rect 11330 1884 11336 1896
rect 11195 1856 11336 1884
rect 11195 1853 11207 1856
rect 11149 1847 11207 1853
rect 11330 1844 11336 1856
rect 11388 1844 11394 1896
rect 11992 1893 12020 1924
rect 12084 1893 12112 1992
rect 12250 1980 12256 1992
rect 12308 1980 12314 2032
rect 11517 1887 11575 1893
rect 11517 1853 11529 1887
rect 11563 1884 11575 1887
rect 11701 1887 11759 1893
rect 11701 1884 11713 1887
rect 11563 1856 11713 1884
rect 11563 1853 11575 1856
rect 11517 1847 11575 1853
rect 11701 1853 11713 1856
rect 11747 1853 11759 1887
rect 11701 1847 11759 1853
rect 11977 1887 12035 1893
rect 11977 1853 11989 1887
rect 12023 1853 12035 1887
rect 11977 1847 12035 1853
rect 12074 1887 12132 1893
rect 12074 1853 12086 1887
rect 12120 1853 12132 1887
rect 12802 1884 12808 1896
rect 12763 1856 12808 1884
rect 12074 1847 12132 1853
rect 12802 1844 12808 1856
rect 12860 1844 12866 1896
rect 12894 1844 12900 1896
rect 12952 1884 12958 1896
rect 13081 1887 13139 1893
rect 13081 1884 13093 1887
rect 12952 1856 13093 1884
rect 12952 1844 12958 1856
rect 13081 1853 13093 1856
rect 13127 1853 13139 1887
rect 13081 1847 13139 1853
rect 11885 1819 11943 1825
rect 11885 1816 11897 1819
rect 11072 1788 11897 1816
rect 11885 1785 11897 1788
rect 11931 1785 11943 1819
rect 11885 1779 11943 1785
rect 12621 1751 12679 1757
rect 12621 1748 12633 1751
rect 10244 1720 12633 1748
rect 12621 1717 12633 1720
rect 12667 1717 12679 1751
rect 12621 1711 12679 1717
rect 1104 1658 13892 1680
rect 1104 1606 8246 1658
rect 8298 1606 8310 1658
rect 8362 1606 8374 1658
rect 8426 1606 8438 1658
rect 8490 1606 13892 1658
rect 1104 1584 13892 1606
rect 2409 1547 2467 1553
rect 2409 1513 2421 1547
rect 2455 1513 2467 1547
rect 2866 1544 2872 1556
rect 2827 1516 2872 1544
rect 2409 1507 2467 1513
rect 2424 1476 2452 1507
rect 2866 1504 2872 1516
rect 2924 1504 2930 1556
rect 6089 1547 6147 1553
rect 6089 1513 6101 1547
rect 6135 1513 6147 1547
rect 6638 1544 6644 1556
rect 6599 1516 6644 1544
rect 6089 1507 6147 1513
rect 6104 1476 6132 1507
rect 6638 1504 6644 1516
rect 6696 1504 6702 1556
rect 6730 1504 6736 1556
rect 6788 1504 6794 1556
rect 8754 1544 8760 1556
rect 8715 1516 8760 1544
rect 8754 1504 8760 1516
rect 8812 1504 8818 1556
rect 9217 1547 9275 1553
rect 9217 1513 9229 1547
rect 9263 1513 9275 1547
rect 9766 1544 9772 1556
rect 9727 1516 9772 1544
rect 9217 1507 9275 1513
rect 6748 1476 6776 1504
rect 2424 1448 5106 1476
rect 6104 1448 6776 1476
rect 1946 1368 1952 1420
rect 2004 1408 2010 1420
rect 2225 1411 2283 1417
rect 2225 1408 2237 1411
rect 2004 1380 2237 1408
rect 2004 1368 2010 1380
rect 2225 1377 2237 1380
rect 2271 1408 2283 1411
rect 2682 1408 2688 1420
rect 2271 1380 2688 1408
rect 2271 1377 2283 1380
rect 2225 1371 2283 1377
rect 2682 1368 2688 1380
rect 2740 1368 2746 1420
rect 3326 1408 3332 1420
rect 3287 1380 3332 1408
rect 3326 1368 3332 1380
rect 3384 1368 3390 1420
rect 3513 1411 3571 1417
rect 3513 1377 3525 1411
rect 3559 1408 3571 1411
rect 3970 1408 3976 1420
rect 3559 1380 3976 1408
rect 3559 1377 3571 1380
rect 3513 1371 3571 1377
rect 3970 1368 3976 1380
rect 4028 1368 4034 1420
rect 4065 1411 4123 1417
rect 4065 1377 4077 1411
rect 4111 1408 4123 1411
rect 4246 1408 4252 1420
rect 4111 1380 4252 1408
rect 4111 1377 4123 1380
rect 4065 1371 4123 1377
rect 4246 1368 4252 1380
rect 4304 1368 4310 1420
rect 6748 1417 6776 1448
rect 7285 1479 7343 1485
rect 7285 1445 7297 1479
rect 7331 1476 7343 1479
rect 7558 1476 7564 1488
rect 7331 1448 7564 1476
rect 7331 1445 7343 1448
rect 7285 1439 7343 1445
rect 7558 1436 7564 1448
rect 7616 1436 7622 1488
rect 9232 1476 9260 1507
rect 9766 1504 9772 1516
rect 9824 1504 9830 1556
rect 11701 1547 11759 1553
rect 11701 1544 11713 1547
rect 9968 1516 11713 1544
rect 9968 1476 9996 1516
rect 11701 1513 11713 1516
rect 11747 1513 11759 1547
rect 11701 1507 11759 1513
rect 11885 1547 11943 1553
rect 11885 1513 11897 1547
rect 11931 1513 11943 1547
rect 11885 1507 11943 1513
rect 12529 1547 12587 1553
rect 12529 1513 12541 1547
rect 12575 1544 12587 1547
rect 12618 1544 12624 1556
rect 12575 1516 12624 1544
rect 12575 1513 12587 1516
rect 12529 1507 12587 1513
rect 11900 1476 11928 1507
rect 12618 1504 12624 1516
rect 12676 1504 12682 1556
rect 8510 1448 9260 1476
rect 9416 1448 9996 1476
rect 10810 1448 11928 1476
rect 9416 1420 9444 1448
rect 6733 1411 6791 1417
rect 6733 1377 6745 1411
rect 6779 1377 6791 1411
rect 9398 1408 9404 1420
rect 9311 1380 9404 1408
rect 6733 1371 6791 1377
rect 9398 1368 9404 1380
rect 9456 1368 9462 1420
rect 11514 1368 11520 1420
rect 11572 1408 11578 1420
rect 11701 1411 11759 1417
rect 11572 1380 11617 1408
rect 11572 1368 11578 1380
rect 11701 1377 11713 1411
rect 11747 1408 11759 1411
rect 12069 1411 12127 1417
rect 12069 1408 12081 1411
rect 11747 1380 12081 1408
rect 11747 1377 11759 1380
rect 11701 1371 11759 1377
rect 12069 1377 12081 1380
rect 12115 1408 12127 1411
rect 12345 1411 12403 1417
rect 12345 1408 12357 1411
rect 12115 1380 12357 1408
rect 12115 1377 12127 1380
rect 12069 1371 12127 1377
rect 12345 1377 12357 1380
rect 12391 1408 12403 1411
rect 12802 1408 12808 1420
rect 12391 1380 12808 1408
rect 12391 1377 12403 1380
rect 12345 1371 12403 1377
rect 12802 1368 12808 1380
rect 12860 1368 12866 1420
rect 4341 1343 4399 1349
rect 4341 1309 4353 1343
rect 4387 1309 4399 1343
rect 4614 1340 4620 1352
rect 4575 1312 4620 1340
rect 4341 1303 4399 1309
rect 3421 1275 3479 1281
rect 3421 1241 3433 1275
rect 3467 1272 3479 1275
rect 4154 1272 4160 1284
rect 3467 1244 4160 1272
rect 3467 1241 3479 1244
rect 3421 1235 3479 1241
rect 4154 1232 4160 1244
rect 4212 1232 4218 1284
rect 4062 1164 4068 1216
rect 4120 1204 4126 1216
rect 4356 1204 4384 1303
rect 4614 1300 4620 1312
rect 4672 1300 4678 1352
rect 6822 1300 6828 1352
rect 6880 1340 6886 1352
rect 7009 1343 7067 1349
rect 7009 1340 7021 1343
rect 6880 1312 7021 1340
rect 6880 1300 6886 1312
rect 7009 1309 7021 1312
rect 7055 1309 7067 1343
rect 7009 1303 7067 1309
rect 11241 1343 11299 1349
rect 11241 1309 11253 1343
rect 11287 1340 11299 1343
rect 12250 1340 12256 1352
rect 11287 1312 12256 1340
rect 11287 1309 11299 1312
rect 11241 1303 11299 1309
rect 12250 1300 12256 1312
rect 12308 1300 12314 1352
rect 6178 1204 6184 1216
rect 4120 1176 6184 1204
rect 4120 1164 4126 1176
rect 6178 1164 6184 1176
rect 6236 1164 6242 1216
rect 1104 1114 13892 1136
rect 1104 1062 4246 1114
rect 4298 1062 4310 1114
rect 4362 1062 4374 1114
rect 4426 1062 4438 1114
rect 4490 1062 12246 1114
rect 12298 1062 12310 1114
rect 12362 1062 12374 1114
rect 12426 1062 12438 1114
rect 12490 1062 13892 1114
rect 1104 1040 13892 1062
<< via1 >>
rect 8246 15750 8298 15802
rect 8310 15750 8362 15802
rect 8374 15750 8426 15802
rect 8438 15750 8490 15802
rect 4620 15648 4672 15700
rect 4988 15580 5040 15632
rect 4896 15512 4948 15564
rect 6552 15512 6604 15564
rect 6828 15555 6880 15564
rect 6828 15521 6837 15555
rect 6837 15521 6871 15555
rect 6871 15521 6880 15555
rect 6828 15512 6880 15521
rect 4804 15444 4856 15496
rect 5816 15444 5868 15496
rect 6460 15444 6512 15496
rect 8760 15512 8812 15564
rect 10232 15555 10284 15564
rect 10232 15521 10241 15555
rect 10241 15521 10275 15555
rect 10275 15521 10284 15555
rect 10232 15512 10284 15521
rect 8024 15487 8076 15496
rect 8024 15453 8033 15487
rect 8033 15453 8067 15487
rect 8067 15453 8076 15487
rect 8024 15444 8076 15453
rect 7012 15376 7064 15428
rect 4068 15351 4120 15360
rect 4068 15317 4077 15351
rect 4077 15317 4111 15351
rect 4111 15317 4120 15351
rect 4068 15308 4120 15317
rect 4620 15308 4672 15360
rect 5448 15351 5500 15360
rect 5448 15317 5457 15351
rect 5457 15317 5491 15351
rect 5491 15317 5500 15351
rect 5448 15308 5500 15317
rect 6644 15351 6696 15360
rect 6644 15317 6653 15351
rect 6653 15317 6687 15351
rect 6687 15317 6696 15351
rect 6644 15308 6696 15317
rect 7288 15351 7340 15360
rect 7288 15317 7297 15351
rect 7297 15317 7331 15351
rect 7331 15317 7340 15351
rect 7288 15308 7340 15317
rect 8576 15308 8628 15360
rect 10140 15351 10192 15360
rect 10140 15317 10149 15351
rect 10149 15317 10183 15351
rect 10183 15317 10192 15351
rect 10140 15308 10192 15317
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 12246 15206 12298 15258
rect 12310 15206 12362 15258
rect 12374 15206 12426 15258
rect 12438 15206 12490 15258
rect 6000 15147 6052 15156
rect 6000 15113 6009 15147
rect 6009 15113 6043 15147
rect 6043 15113 6052 15147
rect 6000 15104 6052 15113
rect 6920 14968 6972 15020
rect 7932 14968 7984 15020
rect 8484 14968 8536 15020
rect 9864 15011 9916 15020
rect 9864 14977 9873 15011
rect 9873 14977 9907 15011
rect 9907 14977 9916 15011
rect 9864 14968 9916 14977
rect 10416 15104 10468 15156
rect 4620 14900 4672 14952
rect 4896 14900 4948 14952
rect 6644 14900 6696 14952
rect 8024 14900 8076 14952
rect 12532 14900 12584 14952
rect 8576 14875 8628 14884
rect 8576 14841 8585 14875
rect 8585 14841 8619 14875
rect 8619 14841 8628 14875
rect 8576 14832 8628 14841
rect 8760 14875 8812 14884
rect 8760 14841 8769 14875
rect 8769 14841 8803 14875
rect 8803 14841 8812 14875
rect 8760 14832 8812 14841
rect 4804 14764 4856 14816
rect 6736 14807 6788 14816
rect 6736 14773 6745 14807
rect 6745 14773 6779 14807
rect 6779 14773 6788 14807
rect 6736 14764 6788 14773
rect 8024 14764 8076 14816
rect 9220 14764 9272 14816
rect 9772 14807 9824 14816
rect 9772 14773 9781 14807
rect 9781 14773 9815 14807
rect 9815 14773 9824 14807
rect 9772 14764 9824 14773
rect 11152 14764 11204 14816
rect 8246 14662 8298 14714
rect 8310 14662 8362 14714
rect 8374 14662 8426 14714
rect 8438 14662 8490 14714
rect 1860 14560 1912 14612
rect 8576 14560 8628 14612
rect 4068 14492 4120 14544
rect 4804 14492 4856 14544
rect 5448 14492 5500 14544
rect 7288 14492 7340 14544
rect 3056 14424 3108 14476
rect 2044 14356 2096 14408
rect 2780 14288 2832 14340
rect 1768 14263 1820 14272
rect 1768 14229 1777 14263
rect 1777 14229 1811 14263
rect 1811 14229 1820 14263
rect 1768 14220 1820 14229
rect 4620 14424 4672 14476
rect 5908 14424 5960 14476
rect 6460 14467 6512 14476
rect 6460 14433 6469 14467
rect 6469 14433 6503 14467
rect 6503 14433 6512 14467
rect 6460 14424 6512 14433
rect 6552 14424 6604 14476
rect 7564 14424 7616 14476
rect 3332 14356 3384 14408
rect 6736 14356 6788 14408
rect 8852 14424 8904 14476
rect 9220 14467 9272 14476
rect 9220 14433 9229 14467
rect 9229 14433 9263 14467
rect 9263 14433 9272 14467
rect 9220 14424 9272 14433
rect 10968 14424 11020 14476
rect 3884 14288 3936 14340
rect 6828 14331 6880 14340
rect 6828 14297 6837 14331
rect 6837 14297 6871 14331
rect 6871 14297 6880 14331
rect 6828 14288 6880 14297
rect 8668 14331 8720 14340
rect 8668 14297 8677 14331
rect 8677 14297 8711 14331
rect 8711 14297 8720 14331
rect 8668 14288 8720 14297
rect 9956 14220 10008 14272
rect 10876 14220 10928 14272
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 12246 14118 12298 14170
rect 12310 14118 12362 14170
rect 12374 14118 12426 14170
rect 12438 14118 12490 14170
rect 5908 14059 5960 14068
rect 5908 14025 5917 14059
rect 5917 14025 5951 14059
rect 5951 14025 5960 14059
rect 5908 14016 5960 14025
rect 8668 14016 8720 14068
rect 4068 13948 4120 14000
rect 3884 13880 3936 13932
rect 6828 13948 6880 14000
rect 8576 13948 8628 14000
rect 9956 13991 10008 14000
rect 9956 13957 9965 13991
rect 9965 13957 9999 13991
rect 9999 13957 10008 13991
rect 9956 13948 10008 13957
rect 10232 13948 10284 14000
rect 11704 13948 11756 14000
rect 7012 13923 7064 13932
rect 1768 13812 1820 13864
rect 3332 13855 3384 13864
rect 3332 13821 3341 13855
rect 3341 13821 3375 13855
rect 3375 13821 3384 13855
rect 3332 13812 3384 13821
rect 4804 13855 4856 13864
rect 4804 13821 4813 13855
rect 4813 13821 4847 13855
rect 4847 13821 4856 13855
rect 4804 13812 4856 13821
rect 7012 13889 7021 13923
rect 7021 13889 7055 13923
rect 7055 13889 7064 13923
rect 7012 13880 7064 13889
rect 9220 13880 9272 13932
rect 10140 13880 10192 13932
rect 10876 13923 10928 13932
rect 10876 13889 10885 13923
rect 10885 13889 10919 13923
rect 10919 13889 10928 13923
rect 10876 13880 10928 13889
rect 12716 13880 12768 13932
rect 5816 13812 5868 13864
rect 7564 13855 7616 13864
rect 7564 13821 7573 13855
rect 7573 13821 7607 13855
rect 7607 13821 7616 13855
rect 7564 13812 7616 13821
rect 8760 13855 8812 13864
rect 8760 13821 8769 13855
rect 8769 13821 8803 13855
rect 8803 13821 8812 13855
rect 8760 13812 8812 13821
rect 10324 13855 10376 13864
rect 10324 13821 10333 13855
rect 10333 13821 10367 13855
rect 10367 13821 10376 13855
rect 10324 13812 10376 13821
rect 10968 13812 11020 13864
rect 12440 13855 12492 13864
rect 12440 13821 12449 13855
rect 12449 13821 12483 13855
rect 12483 13821 12492 13855
rect 12440 13812 12492 13821
rect 13268 13812 13320 13864
rect 2504 13787 2556 13796
rect 2504 13753 2513 13787
rect 2513 13753 2547 13787
rect 2547 13753 2556 13787
rect 2504 13744 2556 13753
rect 2780 13787 2832 13796
rect 2780 13753 2789 13787
rect 2789 13753 2823 13787
rect 2823 13753 2832 13787
rect 11888 13787 11940 13796
rect 2780 13744 2832 13753
rect 11888 13753 11897 13787
rect 11897 13753 11931 13787
rect 11931 13753 11940 13787
rect 11888 13744 11940 13753
rect 5540 13719 5592 13728
rect 5540 13685 5549 13719
rect 5549 13685 5583 13719
rect 5583 13685 5592 13719
rect 5540 13676 5592 13685
rect 11244 13719 11296 13728
rect 11244 13685 11253 13719
rect 11253 13685 11287 13719
rect 11287 13685 11296 13719
rect 11244 13676 11296 13685
rect 11612 13676 11664 13728
rect 12992 13719 13044 13728
rect 12992 13685 13001 13719
rect 13001 13685 13035 13719
rect 13035 13685 13044 13719
rect 12992 13676 13044 13685
rect 8246 13574 8298 13626
rect 8310 13574 8362 13626
rect 8374 13574 8426 13626
rect 8438 13574 8490 13626
rect 2872 13515 2924 13524
rect 2872 13481 2881 13515
rect 2881 13481 2915 13515
rect 2915 13481 2924 13515
rect 2872 13472 2924 13481
rect 3056 13472 3108 13524
rect 2504 13404 2556 13456
rect 4804 13404 4856 13456
rect 6368 13404 6420 13456
rect 6552 13404 6604 13456
rect 1768 13336 1820 13388
rect 3056 13336 3108 13388
rect 2780 13268 2832 13320
rect 4712 13336 4764 13388
rect 5356 13379 5408 13388
rect 5356 13345 5365 13379
rect 5365 13345 5399 13379
rect 5399 13345 5408 13379
rect 5356 13336 5408 13345
rect 5724 13336 5776 13388
rect 5908 13336 5960 13388
rect 6460 13336 6512 13388
rect 8852 13472 8904 13524
rect 9312 13472 9364 13524
rect 8576 13404 8628 13456
rect 8760 13404 8812 13456
rect 10232 13447 10284 13456
rect 10232 13413 10241 13447
rect 10241 13413 10275 13447
rect 10275 13413 10284 13447
rect 10232 13404 10284 13413
rect 10968 13404 11020 13456
rect 12440 13404 12492 13456
rect 13176 13404 13228 13456
rect 5172 13268 5224 13320
rect 7656 13336 7708 13388
rect 8116 13336 8168 13388
rect 9496 13336 9548 13388
rect 9680 13336 9732 13388
rect 10324 13336 10376 13388
rect 7932 13268 7984 13320
rect 8852 13268 8904 13320
rect 10416 13268 10468 13320
rect 7380 13200 7432 13252
rect 11612 13336 11664 13388
rect 12716 13379 12768 13388
rect 12716 13345 12725 13379
rect 12725 13345 12759 13379
rect 12759 13345 12768 13379
rect 12716 13336 12768 13345
rect 13360 13379 13412 13388
rect 13360 13345 13369 13379
rect 13369 13345 13403 13379
rect 13403 13345 13412 13379
rect 13360 13336 13412 13345
rect 11336 13200 11388 13252
rect 2964 13132 3016 13184
rect 5080 13175 5132 13184
rect 5080 13141 5089 13175
rect 5089 13141 5123 13175
rect 5123 13141 5132 13175
rect 5080 13132 5132 13141
rect 6828 13132 6880 13184
rect 10968 13132 11020 13184
rect 13084 13132 13136 13184
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 12246 13030 12298 13082
rect 12310 13030 12362 13082
rect 12374 13030 12426 13082
rect 12438 13030 12490 13082
rect 2044 12860 2096 12912
rect 5080 12928 5132 12980
rect 7564 12928 7616 12980
rect 8024 12928 8076 12980
rect 8944 12928 8996 12980
rect 9680 12928 9732 12980
rect 3056 12860 3108 12912
rect 3240 12860 3292 12912
rect 4344 12860 4396 12912
rect 6552 12860 6604 12912
rect 2964 12835 3016 12844
rect 2964 12801 2973 12835
rect 2973 12801 3007 12835
rect 3007 12801 3016 12835
rect 2964 12792 3016 12801
rect 4712 12792 4764 12844
rect 5816 12792 5868 12844
rect 8852 12835 8904 12844
rect 3148 12724 3200 12776
rect 1676 12631 1728 12640
rect 1676 12597 1685 12631
rect 1685 12597 1719 12631
rect 1719 12597 1728 12631
rect 1676 12588 1728 12597
rect 2136 12631 2188 12640
rect 2136 12597 2145 12631
rect 2145 12597 2179 12631
rect 2179 12597 2188 12631
rect 2136 12588 2188 12597
rect 4804 12656 4856 12708
rect 5356 12656 5408 12708
rect 6276 12656 6328 12708
rect 6920 12699 6972 12708
rect 6920 12665 6929 12699
rect 6929 12665 6963 12699
rect 6963 12665 6972 12699
rect 6920 12656 6972 12665
rect 8852 12801 8861 12835
rect 8861 12801 8895 12835
rect 8895 12801 8904 12835
rect 8852 12792 8904 12801
rect 7472 12724 7524 12776
rect 7748 12724 7800 12776
rect 10876 12860 10928 12912
rect 9864 12792 9916 12844
rect 10232 12835 10284 12844
rect 10232 12801 10241 12835
rect 10241 12801 10275 12835
rect 10275 12801 10284 12835
rect 10232 12792 10284 12801
rect 10416 12835 10468 12844
rect 10416 12801 10425 12835
rect 10425 12801 10459 12835
rect 10459 12801 10468 12835
rect 10416 12792 10468 12801
rect 11244 12792 11296 12844
rect 11796 12724 11848 12776
rect 13176 12767 13228 12776
rect 13176 12733 13185 12767
rect 13185 12733 13219 12767
rect 13219 12733 13228 12767
rect 13176 12724 13228 12733
rect 7932 12656 7984 12708
rect 8024 12656 8076 12708
rect 8668 12656 8720 12708
rect 8852 12656 8904 12708
rect 11888 12656 11940 12708
rect 6000 12588 6052 12640
rect 7012 12631 7064 12640
rect 7012 12597 7021 12631
rect 7021 12597 7055 12631
rect 7055 12597 7064 12631
rect 7012 12588 7064 12597
rect 7380 12631 7432 12640
rect 7380 12597 7389 12631
rect 7389 12597 7423 12631
rect 7423 12597 7432 12631
rect 7380 12588 7432 12597
rect 8576 12588 8628 12640
rect 9220 12588 9272 12640
rect 8246 12486 8298 12538
rect 8310 12486 8362 12538
rect 8374 12486 8426 12538
rect 8438 12486 8490 12538
rect 4344 12427 4396 12436
rect 4344 12393 4353 12427
rect 4353 12393 4387 12427
rect 4387 12393 4396 12427
rect 4344 12384 4396 12393
rect 5540 12384 5592 12436
rect 7012 12384 7064 12436
rect 7196 12384 7248 12436
rect 3056 12359 3108 12368
rect 3056 12325 3065 12359
rect 3065 12325 3099 12359
rect 3099 12325 3108 12359
rect 3056 12316 3108 12325
rect 4804 12316 4856 12368
rect 5264 12316 5316 12368
rect 9128 12384 9180 12436
rect 9312 12427 9364 12436
rect 9312 12393 9321 12427
rect 9321 12393 9355 12427
rect 9355 12393 9364 12427
rect 9312 12384 9364 12393
rect 10324 12384 10376 12436
rect 11428 12384 11480 12436
rect 13176 12384 13228 12436
rect 2136 12248 2188 12300
rect 2780 12291 2832 12300
rect 2780 12257 2789 12291
rect 2789 12257 2823 12291
rect 2823 12257 2832 12291
rect 2780 12248 2832 12257
rect 4068 12248 4120 12300
rect 5172 12291 5224 12300
rect 5172 12257 5181 12291
rect 5181 12257 5215 12291
rect 5215 12257 5224 12291
rect 5172 12248 5224 12257
rect 2044 12180 2096 12232
rect 5448 12291 5500 12300
rect 5448 12257 5457 12291
rect 5457 12257 5491 12291
rect 5491 12257 5500 12291
rect 5448 12248 5500 12257
rect 7564 12316 7616 12368
rect 9496 12316 9548 12368
rect 10232 12316 10284 12368
rect 11704 12359 11756 12368
rect 7380 12248 7432 12300
rect 7748 12291 7800 12300
rect 7748 12257 7757 12291
rect 7757 12257 7791 12291
rect 7791 12257 7800 12291
rect 7748 12248 7800 12257
rect 8024 12248 8076 12300
rect 8484 12291 8536 12300
rect 8484 12257 8493 12291
rect 8493 12257 8527 12291
rect 8527 12257 8536 12291
rect 8484 12248 8536 12257
rect 8760 12248 8812 12300
rect 10140 12248 10192 12300
rect 11704 12325 11713 12359
rect 11713 12325 11747 12359
rect 11747 12325 11756 12359
rect 11704 12316 11756 12325
rect 10600 12248 10652 12300
rect 11336 12248 11388 12300
rect 11612 12291 11664 12300
rect 11612 12257 11621 12291
rect 11621 12257 11655 12291
rect 11655 12257 11664 12291
rect 11612 12248 11664 12257
rect 13176 12291 13228 12300
rect 13176 12257 13185 12291
rect 13185 12257 13219 12291
rect 13219 12257 13228 12291
rect 13176 12248 13228 12257
rect 3148 12112 3200 12164
rect 6828 12180 6880 12232
rect 8116 12180 8168 12232
rect 8392 12180 8444 12232
rect 4896 12112 4948 12164
rect 6092 12112 6144 12164
rect 3792 12044 3844 12096
rect 5172 12044 5224 12096
rect 5632 12044 5684 12096
rect 7288 12112 7340 12164
rect 12072 12180 12124 12232
rect 10416 12112 10468 12164
rect 12808 12112 12860 12164
rect 6368 12044 6420 12096
rect 6920 12044 6972 12096
rect 7012 12044 7064 12096
rect 8484 12087 8536 12096
rect 8484 12053 8493 12087
rect 8493 12053 8527 12087
rect 8527 12053 8536 12087
rect 8484 12044 8536 12053
rect 9312 12044 9364 12096
rect 11980 12087 12032 12096
rect 11980 12053 11989 12087
rect 11989 12053 12023 12087
rect 12023 12053 12032 12087
rect 11980 12044 12032 12053
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 12246 11942 12298 11994
rect 12310 11942 12362 11994
rect 12374 11942 12426 11994
rect 12438 11942 12490 11994
rect 6000 11883 6052 11892
rect 6000 11849 6009 11883
rect 6009 11849 6043 11883
rect 6043 11849 6052 11883
rect 6000 11840 6052 11849
rect 6552 11883 6604 11892
rect 6552 11849 6561 11883
rect 6561 11849 6595 11883
rect 6595 11849 6604 11883
rect 6552 11840 6604 11849
rect 5080 11815 5132 11824
rect 5080 11781 5089 11815
rect 5089 11781 5123 11815
rect 5123 11781 5132 11815
rect 5080 11772 5132 11781
rect 6736 11772 6788 11824
rect 480 11704 532 11756
rect 2044 11636 2096 11688
rect 3148 11679 3200 11688
rect 3148 11645 3157 11679
rect 3157 11645 3191 11679
rect 3191 11645 3200 11679
rect 3148 11636 3200 11645
rect 3424 11679 3476 11688
rect 3424 11645 3433 11679
rect 3433 11645 3467 11679
rect 3467 11645 3476 11679
rect 3424 11636 3476 11645
rect 1768 11543 1820 11552
rect 1768 11509 1777 11543
rect 1777 11509 1811 11543
rect 1811 11509 1820 11543
rect 1768 11500 1820 11509
rect 2780 11611 2832 11620
rect 2780 11577 2789 11611
rect 2789 11577 2823 11611
rect 2823 11577 2832 11611
rect 2780 11568 2832 11577
rect 3332 11568 3384 11620
rect 5540 11704 5592 11756
rect 6092 11704 6144 11756
rect 8484 11840 8536 11892
rect 10140 11840 10192 11892
rect 8576 11772 8628 11824
rect 9220 11772 9272 11824
rect 11796 11840 11848 11892
rect 13176 11815 13228 11824
rect 13176 11781 13185 11815
rect 13185 11781 13219 11815
rect 13219 11781 13228 11815
rect 13176 11772 13228 11781
rect 7288 11704 7340 11756
rect 8392 11747 8444 11756
rect 8392 11713 8401 11747
rect 8401 11713 8435 11747
rect 8435 11713 8444 11747
rect 8392 11704 8444 11713
rect 3976 11636 4028 11688
rect 6460 11636 6512 11688
rect 7380 11636 7432 11688
rect 8024 11679 8076 11688
rect 8024 11645 8033 11679
rect 8033 11645 8067 11679
rect 8067 11645 8076 11679
rect 8024 11636 8076 11645
rect 8852 11704 8904 11756
rect 9128 11704 9180 11756
rect 9680 11704 9732 11756
rect 10508 11747 10560 11756
rect 10508 11713 10517 11747
rect 10517 11713 10551 11747
rect 10551 11713 10560 11747
rect 10508 11704 10560 11713
rect 12808 11704 12860 11756
rect 13268 11747 13320 11756
rect 13268 11713 13277 11747
rect 13277 11713 13311 11747
rect 13311 11713 13320 11747
rect 13268 11704 13320 11713
rect 8668 11679 8720 11688
rect 8668 11645 8677 11679
rect 8677 11645 8711 11679
rect 8711 11645 8720 11679
rect 8668 11636 8720 11645
rect 9312 11679 9364 11688
rect 9312 11645 9321 11679
rect 9321 11645 9355 11679
rect 9355 11645 9364 11679
rect 9312 11636 9364 11645
rect 10968 11679 11020 11688
rect 4068 11568 4120 11620
rect 5264 11611 5316 11620
rect 5264 11577 5273 11611
rect 5273 11577 5307 11611
rect 5307 11577 5316 11611
rect 5264 11568 5316 11577
rect 5632 11611 5684 11620
rect 5632 11577 5641 11611
rect 5641 11577 5675 11611
rect 5675 11577 5684 11611
rect 5632 11568 5684 11577
rect 6368 11568 6420 11620
rect 8116 11568 8168 11620
rect 9404 11568 9456 11620
rect 10232 11568 10284 11620
rect 10968 11645 10977 11679
rect 10977 11645 11011 11679
rect 11011 11645 11020 11679
rect 10968 11636 11020 11645
rect 11796 11636 11848 11688
rect 11980 11636 12032 11688
rect 4712 11500 4764 11552
rect 5356 11543 5408 11552
rect 5356 11509 5365 11543
rect 5365 11509 5399 11543
rect 5399 11509 5408 11543
rect 5356 11500 5408 11509
rect 5724 11500 5776 11552
rect 5908 11500 5960 11552
rect 8668 11500 8720 11552
rect 9864 11500 9916 11552
rect 11888 11500 11940 11552
rect 8246 11398 8298 11450
rect 8310 11398 8362 11450
rect 8374 11398 8426 11450
rect 8438 11398 8490 11450
rect 3424 11296 3476 11348
rect 1768 11203 1820 11212
rect 1768 11169 1777 11203
rect 1777 11169 1811 11203
rect 1811 11169 1820 11203
rect 1768 11160 1820 11169
rect 2412 11203 2464 11212
rect 2412 11169 2421 11203
rect 2421 11169 2455 11203
rect 2455 11169 2464 11203
rect 2412 11160 2464 11169
rect 2688 11203 2740 11212
rect 2688 11169 2697 11203
rect 2697 11169 2731 11203
rect 2731 11169 2740 11203
rect 2688 11160 2740 11169
rect 3792 11228 3844 11280
rect 3976 11271 4028 11280
rect 3976 11237 3985 11271
rect 3985 11237 4019 11271
rect 4019 11237 4028 11271
rect 3976 11228 4028 11237
rect 8024 11339 8076 11348
rect 8024 11305 8033 11339
rect 8033 11305 8067 11339
rect 8067 11305 8076 11339
rect 8024 11296 8076 11305
rect 9772 11296 9824 11348
rect 10508 11296 10560 11348
rect 5908 11228 5960 11280
rect 7840 11228 7892 11280
rect 9036 11228 9088 11280
rect 10048 11228 10100 11280
rect 10968 11271 11020 11280
rect 10968 11237 10977 11271
rect 10977 11237 11011 11271
rect 11011 11237 11020 11271
rect 10968 11228 11020 11237
rect 13176 11228 13228 11280
rect 5080 11160 5132 11212
rect 5172 11203 5224 11212
rect 5172 11169 5181 11203
rect 5181 11169 5215 11203
rect 5215 11169 5224 11203
rect 5448 11203 5500 11212
rect 5172 11160 5224 11169
rect 5448 11169 5457 11203
rect 5457 11169 5491 11203
rect 5491 11169 5500 11203
rect 5448 11160 5500 11169
rect 6000 11203 6052 11212
rect 6000 11169 6009 11203
rect 6009 11169 6043 11203
rect 6043 11169 6052 11203
rect 6000 11160 6052 11169
rect 6460 11203 6512 11212
rect 6460 11169 6469 11203
rect 6469 11169 6503 11203
rect 6503 11169 6512 11203
rect 6460 11160 6512 11169
rect 6736 11203 6788 11212
rect 6736 11169 6745 11203
rect 6745 11169 6779 11203
rect 6779 11169 6788 11203
rect 6736 11160 6788 11169
rect 7012 11203 7064 11212
rect 7012 11169 7021 11203
rect 7021 11169 7055 11203
rect 7055 11169 7064 11203
rect 7012 11160 7064 11169
rect 7196 11203 7248 11212
rect 7196 11169 7205 11203
rect 7205 11169 7239 11203
rect 7239 11169 7248 11203
rect 7196 11160 7248 11169
rect 7932 11160 7984 11212
rect 2964 11135 3016 11144
rect 2964 11101 2973 11135
rect 2973 11101 3007 11135
rect 3007 11101 3016 11135
rect 2964 11092 3016 11101
rect 6092 11092 6144 11144
rect 6920 11135 6972 11144
rect 6920 11101 6929 11135
rect 6929 11101 6963 11135
rect 6963 11101 6972 11135
rect 6920 11092 6972 11101
rect 8668 11160 8720 11212
rect 9956 11203 10008 11212
rect 9956 11169 9965 11203
rect 9965 11169 9999 11203
rect 9999 11169 10008 11203
rect 9956 11160 10008 11169
rect 8852 11092 8904 11144
rect 10784 11160 10836 11212
rect 11980 11160 12032 11212
rect 13268 11203 13320 11212
rect 13268 11169 13277 11203
rect 13277 11169 13311 11203
rect 13311 11169 13320 11203
rect 13268 11160 13320 11169
rect 2412 11024 2464 11076
rect 4804 11024 4856 11076
rect 5724 11024 5776 11076
rect 6828 11067 6880 11076
rect 6828 11033 6837 11067
rect 6837 11033 6871 11067
rect 6871 11033 6880 11067
rect 6828 11024 6880 11033
rect 9128 11024 9180 11076
rect 10600 11092 10652 11144
rect 5816 10956 5868 11008
rect 9220 10956 9272 11008
rect 9864 10956 9916 11008
rect 10416 10956 10468 11008
rect 10600 10999 10652 11008
rect 10600 10965 10609 10999
rect 10609 10965 10643 10999
rect 10643 10965 10652 10999
rect 10600 10956 10652 10965
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 12246 10854 12298 10906
rect 12310 10854 12362 10906
rect 12374 10854 12426 10906
rect 12438 10854 12490 10906
rect 2964 10752 3016 10804
rect 4620 10727 4672 10736
rect 4620 10693 4629 10727
rect 4629 10693 4663 10727
rect 4663 10693 4672 10727
rect 4620 10684 4672 10693
rect 2412 10616 2464 10668
rect 5264 10616 5316 10668
rect 6000 10752 6052 10804
rect 6828 10795 6880 10804
rect 6828 10761 6837 10795
rect 6837 10761 6871 10795
rect 6871 10761 6880 10795
rect 6828 10752 6880 10761
rect 7840 10752 7892 10804
rect 9588 10752 9640 10804
rect 11152 10752 11204 10804
rect 12624 10684 12676 10736
rect 7012 10659 7064 10668
rect 1860 10591 1912 10600
rect 1860 10557 1869 10591
rect 1869 10557 1903 10591
rect 1903 10557 1912 10591
rect 1860 10548 1912 10557
rect 2688 10591 2740 10600
rect 2688 10557 2697 10591
rect 2697 10557 2731 10591
rect 2731 10557 2740 10591
rect 2688 10548 2740 10557
rect 2780 10548 2832 10600
rect 5448 10591 5500 10600
rect 2964 10480 3016 10532
rect 4068 10480 4120 10532
rect 5448 10557 5457 10591
rect 5457 10557 5491 10591
rect 5491 10557 5500 10591
rect 5448 10548 5500 10557
rect 7012 10625 7021 10659
rect 7021 10625 7055 10659
rect 7055 10625 7064 10659
rect 7012 10616 7064 10625
rect 7472 10616 7524 10668
rect 9956 10616 10008 10668
rect 5356 10480 5408 10532
rect 5908 10548 5960 10600
rect 6736 10480 6788 10532
rect 7288 10548 7340 10600
rect 8852 10591 8904 10600
rect 7840 10523 7892 10532
rect 7840 10489 7849 10523
rect 7849 10489 7883 10523
rect 7883 10489 7892 10523
rect 7840 10480 7892 10489
rect 7932 10480 7984 10532
rect 8852 10557 8861 10591
rect 8861 10557 8895 10591
rect 8895 10557 8904 10591
rect 8852 10548 8904 10557
rect 9312 10591 9364 10600
rect 9312 10557 9321 10591
rect 9321 10557 9355 10591
rect 9355 10557 9364 10591
rect 9312 10548 9364 10557
rect 9864 10548 9916 10600
rect 10232 10616 10284 10668
rect 10508 10616 10560 10668
rect 10600 10616 10652 10668
rect 10968 10616 11020 10668
rect 11152 10548 11204 10600
rect 11796 10548 11848 10600
rect 12348 10591 12400 10600
rect 12348 10557 12357 10591
rect 12357 10557 12391 10591
rect 12391 10557 12400 10591
rect 12348 10548 12400 10557
rect 12992 10591 13044 10600
rect 12992 10557 13001 10591
rect 13001 10557 13035 10591
rect 13035 10557 13044 10591
rect 12992 10548 13044 10557
rect 13268 10591 13320 10600
rect 13268 10557 13277 10591
rect 13277 10557 13311 10591
rect 13311 10557 13320 10591
rect 13268 10548 13320 10557
rect 9220 10480 9272 10532
rect 3976 10412 4028 10464
rect 7104 10412 7156 10464
rect 7748 10412 7800 10464
rect 9956 10412 10008 10464
rect 10416 10412 10468 10464
rect 11428 10480 11480 10532
rect 11152 10412 11204 10464
rect 12532 10412 12584 10464
rect 8246 10310 8298 10362
rect 8310 10310 8362 10362
rect 8374 10310 8426 10362
rect 8438 10310 8490 10362
rect 5172 10208 5224 10260
rect 5448 10208 5500 10260
rect 2964 10183 3016 10192
rect 2964 10149 2973 10183
rect 2973 10149 3007 10183
rect 3007 10149 3016 10183
rect 2964 10140 3016 10149
rect 1400 10115 1452 10124
rect 1400 10081 1409 10115
rect 1409 10081 1443 10115
rect 1443 10081 1452 10115
rect 1400 10072 1452 10081
rect 1860 10072 1912 10124
rect 2688 10115 2740 10124
rect 2688 10081 2697 10115
rect 2697 10081 2731 10115
rect 2731 10081 2740 10115
rect 2688 10072 2740 10081
rect 4620 10140 4672 10192
rect 4988 10140 5040 10192
rect 5816 10140 5868 10192
rect 3424 10072 3476 10124
rect 4896 10072 4948 10124
rect 5172 10115 5224 10124
rect 5172 10081 5181 10115
rect 5181 10081 5215 10115
rect 5215 10081 5224 10115
rect 5172 10072 5224 10081
rect 5356 10072 5408 10124
rect 5908 10072 5960 10124
rect 6552 10115 6604 10124
rect 6552 10081 6561 10115
rect 6561 10081 6595 10115
rect 6595 10081 6604 10115
rect 6552 10072 6604 10081
rect 6736 10208 6788 10260
rect 6920 10115 6972 10124
rect 6920 10081 6929 10115
rect 6929 10081 6963 10115
rect 6963 10081 6972 10115
rect 6920 10072 6972 10081
rect 5632 10004 5684 10056
rect 6368 10004 6420 10056
rect 6644 10004 6696 10056
rect 8760 10208 8812 10260
rect 10140 10208 10192 10260
rect 11704 10208 11756 10260
rect 10232 10140 10284 10192
rect 7748 10072 7800 10124
rect 8024 10115 8076 10124
rect 8024 10081 8033 10115
rect 8033 10081 8067 10115
rect 8067 10081 8076 10115
rect 8024 10072 8076 10081
rect 8116 10072 8168 10124
rect 8576 10115 8628 10124
rect 8576 10081 8585 10115
rect 8585 10081 8619 10115
rect 8619 10081 8628 10115
rect 8576 10072 8628 10081
rect 8668 10072 8720 10124
rect 9312 10115 9364 10124
rect 9312 10081 9321 10115
rect 9321 10081 9355 10115
rect 9355 10081 9364 10115
rect 9312 10072 9364 10081
rect 9496 10115 9548 10124
rect 9496 10081 9505 10115
rect 9505 10081 9539 10115
rect 9539 10081 9548 10115
rect 9496 10072 9548 10081
rect 9772 10072 9824 10124
rect 10600 10140 10652 10192
rect 12716 10140 12768 10192
rect 13084 10183 13136 10192
rect 13084 10149 13093 10183
rect 13093 10149 13127 10183
rect 13127 10149 13136 10183
rect 13084 10140 13136 10149
rect 12992 10115 13044 10124
rect 12992 10081 13001 10115
rect 13001 10081 13035 10115
rect 13035 10081 13044 10115
rect 12992 10072 13044 10081
rect 3976 9979 4028 9988
rect 3976 9945 3985 9979
rect 3985 9945 4019 9979
rect 4019 9945 4028 9979
rect 3976 9936 4028 9945
rect 4068 9936 4120 9988
rect 8760 10004 8812 10056
rect 10692 10047 10744 10056
rect 10692 10013 10701 10047
rect 10701 10013 10735 10047
rect 10735 10013 10744 10047
rect 10692 10004 10744 10013
rect 12072 10004 12124 10056
rect 12348 10004 12400 10056
rect 4620 9868 4672 9920
rect 4896 9911 4948 9920
rect 4896 9877 4905 9911
rect 4905 9877 4939 9911
rect 4939 9877 4948 9911
rect 4896 9868 4948 9877
rect 5448 9868 5500 9920
rect 5816 9868 5868 9920
rect 6092 9868 6144 9920
rect 7840 9936 7892 9988
rect 8576 9979 8628 9988
rect 8576 9945 8585 9979
rect 8585 9945 8619 9979
rect 8619 9945 8628 9979
rect 8576 9936 8628 9945
rect 7380 9868 7432 9920
rect 11980 9868 12032 9920
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 12246 9766 12298 9818
rect 12310 9766 12362 9818
rect 12374 9766 12426 9818
rect 12438 9766 12490 9818
rect 1400 9707 1452 9716
rect 1400 9673 1409 9707
rect 1409 9673 1443 9707
rect 1443 9673 1452 9707
rect 1400 9664 1452 9673
rect 3332 9707 3384 9716
rect 3332 9673 3341 9707
rect 3341 9673 3375 9707
rect 3375 9673 3384 9707
rect 3332 9664 3384 9673
rect 5540 9707 5592 9716
rect 5540 9673 5549 9707
rect 5549 9673 5583 9707
rect 5583 9673 5592 9707
rect 5540 9664 5592 9673
rect 5724 9707 5776 9716
rect 5724 9673 5733 9707
rect 5733 9673 5767 9707
rect 5767 9673 5776 9707
rect 5724 9664 5776 9673
rect 7012 9664 7064 9716
rect 4896 9596 4948 9648
rect 6828 9596 6880 9648
rect 9220 9664 9272 9716
rect 10416 9664 10468 9716
rect 10692 9664 10744 9716
rect 12072 9664 12124 9716
rect 8944 9639 8996 9648
rect 2044 9571 2096 9580
rect 2044 9537 2053 9571
rect 2053 9537 2087 9571
rect 2087 9537 2096 9571
rect 2044 9528 2096 9537
rect 5632 9528 5684 9580
rect 8944 9605 8953 9639
rect 8953 9605 8987 9639
rect 8987 9605 8996 9639
rect 8944 9596 8996 9605
rect 2872 9460 2924 9512
rect 3240 9503 3292 9512
rect 3240 9469 3249 9503
rect 3249 9469 3283 9503
rect 3283 9469 3292 9503
rect 3240 9460 3292 9469
rect 3516 9503 3568 9512
rect 3516 9469 3525 9503
rect 3525 9469 3559 9503
rect 3559 9469 3568 9503
rect 3516 9460 3568 9469
rect 4620 9503 4672 9512
rect 4620 9469 4629 9503
rect 4629 9469 4663 9503
rect 4663 9469 4672 9503
rect 4620 9460 4672 9469
rect 5264 9460 5316 9512
rect 3608 9392 3660 9444
rect 5632 9392 5684 9444
rect 5816 9392 5868 9444
rect 7932 9460 7984 9512
rect 9128 9596 9180 9648
rect 10784 9528 10836 9580
rect 12808 9571 12860 9580
rect 12808 9537 12817 9571
rect 12817 9537 12851 9571
rect 12851 9537 12860 9571
rect 12808 9528 12860 9537
rect 7380 9435 7432 9444
rect 1492 9324 1544 9376
rect 2780 9324 2832 9376
rect 5448 9324 5500 9376
rect 7380 9401 7389 9435
rect 7389 9401 7423 9435
rect 7423 9401 7432 9435
rect 7380 9392 7432 9401
rect 7472 9392 7524 9444
rect 8116 9392 8168 9444
rect 8668 9392 8720 9444
rect 7012 9324 7064 9376
rect 7932 9324 7984 9376
rect 9220 9503 9272 9512
rect 9220 9469 9228 9503
rect 9228 9469 9262 9503
rect 9262 9469 9272 9503
rect 9496 9503 9548 9512
rect 9220 9460 9272 9469
rect 9496 9469 9505 9503
rect 9505 9469 9539 9503
rect 9539 9469 9548 9503
rect 9496 9460 9548 9469
rect 9312 9435 9364 9444
rect 9312 9401 9321 9435
rect 9321 9401 9355 9435
rect 9355 9401 9364 9435
rect 9312 9392 9364 9401
rect 10968 9460 11020 9512
rect 9864 9324 9916 9376
rect 10416 9324 10468 9376
rect 11152 9392 11204 9444
rect 11980 9460 12032 9512
rect 12624 9503 12676 9512
rect 12624 9469 12633 9503
rect 12633 9469 12667 9503
rect 12667 9469 12676 9503
rect 12624 9460 12676 9469
rect 10784 9324 10836 9376
rect 13820 9324 13872 9376
rect 8246 9222 8298 9274
rect 8310 9222 8362 9274
rect 8374 9222 8426 9274
rect 8438 9222 8490 9274
rect 2136 8984 2188 9036
rect 2320 9027 2372 9036
rect 2320 8993 2329 9027
rect 2329 8993 2363 9027
rect 2363 8993 2372 9027
rect 2320 8984 2372 8993
rect 3056 9052 3108 9104
rect 3332 9052 3384 9104
rect 4988 9120 5040 9172
rect 5172 9120 5224 9172
rect 5540 9120 5592 9172
rect 6828 9120 6880 9172
rect 5264 9052 5316 9104
rect 6092 9052 6144 9104
rect 7472 9052 7524 9104
rect 3332 8959 3384 8968
rect 3332 8925 3341 8959
rect 3341 8925 3375 8959
rect 3375 8925 3384 8959
rect 3332 8916 3384 8925
rect 4712 8984 4764 9036
rect 4896 9027 4948 9036
rect 4896 8993 4905 9027
rect 4905 8993 4939 9027
rect 4939 8993 4948 9027
rect 4896 8984 4948 8993
rect 5172 9027 5224 9036
rect 4620 8916 4672 8968
rect 5172 8993 5181 9027
rect 5181 8993 5215 9027
rect 5215 8993 5224 9027
rect 5172 8984 5224 8993
rect 7564 8984 7616 9036
rect 8760 9052 8812 9104
rect 9496 9120 9548 9172
rect 9588 9120 9640 9172
rect 10784 9163 10836 9172
rect 10784 9129 10793 9163
rect 10793 9129 10827 9163
rect 10827 9129 10836 9163
rect 10784 9120 10836 9129
rect 12716 9163 12768 9172
rect 8576 8984 8628 9036
rect 9220 8984 9272 9036
rect 9404 9052 9456 9104
rect 10416 9095 10468 9104
rect 10416 9061 10425 9095
rect 10425 9061 10459 9095
rect 10459 9061 10468 9095
rect 10416 9052 10468 9061
rect 2872 8891 2924 8900
rect 2872 8857 2881 8891
rect 2881 8857 2915 8891
rect 2915 8857 2924 8891
rect 2872 8848 2924 8857
rect 5448 8848 5500 8900
rect 1768 8780 1820 8832
rect 5724 8848 5776 8900
rect 7472 8916 7524 8968
rect 7840 8848 7892 8900
rect 8208 8959 8260 8968
rect 8208 8925 8217 8959
rect 8217 8925 8251 8959
rect 8251 8925 8260 8959
rect 8208 8916 8260 8925
rect 10600 9027 10652 9036
rect 10600 8993 10614 9027
rect 10614 8993 10648 9027
rect 10648 8993 10652 9027
rect 10600 8984 10652 8993
rect 11152 9027 11204 9036
rect 11152 8993 11161 9027
rect 11161 8993 11195 9027
rect 11195 8993 11204 9027
rect 11336 9027 11388 9036
rect 11152 8984 11204 8993
rect 11336 8993 11345 9027
rect 11345 8993 11379 9027
rect 11379 8993 11388 9027
rect 11336 8984 11388 8993
rect 11796 9027 11848 9036
rect 11796 8993 11805 9027
rect 11805 8993 11839 9027
rect 11839 8993 11848 9027
rect 11796 8984 11848 8993
rect 12716 9129 12725 9163
rect 12725 9129 12759 9163
rect 12759 9129 12768 9163
rect 12716 9120 12768 9129
rect 12900 9027 12952 9036
rect 12900 8993 12909 9027
rect 12909 8993 12943 9027
rect 12943 8993 12952 9027
rect 12900 8984 12952 8993
rect 8760 8848 8812 8900
rect 8944 8848 8996 8900
rect 11152 8848 11204 8900
rect 11980 8848 12032 8900
rect 6736 8780 6788 8832
rect 7104 8780 7156 8832
rect 8116 8780 8168 8832
rect 9128 8780 9180 8832
rect 9496 8780 9548 8832
rect 9680 8780 9732 8832
rect 9864 8780 9916 8832
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 12246 8678 12298 8730
rect 12310 8678 12362 8730
rect 12374 8678 12426 8730
rect 12438 8678 12490 8730
rect 5356 8619 5408 8628
rect 5356 8585 5365 8619
rect 5365 8585 5399 8619
rect 5399 8585 5408 8619
rect 5356 8576 5408 8585
rect 6092 8619 6144 8628
rect 6092 8585 6101 8619
rect 6101 8585 6135 8619
rect 6135 8585 6144 8619
rect 6092 8576 6144 8585
rect 7104 8619 7156 8628
rect 7104 8585 7113 8619
rect 7113 8585 7147 8619
rect 7147 8585 7156 8619
rect 7104 8576 7156 8585
rect 8668 8619 8720 8628
rect 8668 8585 8677 8619
rect 8677 8585 8711 8619
rect 8711 8585 8720 8619
rect 8668 8576 8720 8585
rect 8760 8576 8812 8628
rect 11336 8576 11388 8628
rect 3332 8508 3384 8560
rect 7932 8508 7984 8560
rect 8208 8551 8260 8560
rect 8208 8517 8217 8551
rect 8217 8517 8251 8551
rect 8251 8517 8260 8551
rect 8208 8508 8260 8517
rect 9220 8508 9272 8560
rect 2044 8483 2096 8492
rect 2044 8449 2053 8483
rect 2053 8449 2087 8483
rect 2087 8449 2096 8483
rect 2044 8440 2096 8449
rect 1768 8415 1820 8424
rect 1768 8381 1777 8415
rect 1777 8381 1811 8415
rect 1811 8381 1820 8415
rect 1768 8372 1820 8381
rect 2872 8372 2924 8424
rect 6184 8440 6236 8492
rect 7012 8483 7064 8492
rect 7012 8449 7021 8483
rect 7021 8449 7055 8483
rect 7055 8449 7064 8483
rect 7012 8440 7064 8449
rect 3608 8415 3660 8424
rect 3608 8381 3617 8415
rect 3617 8381 3651 8415
rect 3651 8381 3660 8415
rect 3608 8372 3660 8381
rect 5816 8372 5868 8424
rect 6828 8415 6880 8424
rect 6828 8381 6837 8415
rect 6837 8381 6871 8415
rect 6871 8381 6880 8415
rect 6828 8372 6880 8381
rect 1860 8347 1912 8356
rect 1860 8313 1869 8347
rect 1869 8313 1903 8347
rect 1903 8313 1912 8347
rect 1860 8304 1912 8313
rect 2412 8347 2464 8356
rect 2412 8313 2421 8347
rect 2421 8313 2455 8347
rect 2455 8313 2464 8347
rect 2412 8304 2464 8313
rect 4160 8304 4212 8356
rect 5632 8304 5684 8356
rect 7564 8372 7616 8424
rect 7748 8372 7800 8424
rect 1400 8279 1452 8288
rect 1400 8245 1409 8279
rect 1409 8245 1443 8279
rect 1443 8245 1452 8279
rect 1400 8236 1452 8245
rect 4896 8236 4948 8288
rect 7288 8304 7340 8356
rect 8116 8304 8168 8356
rect 8760 8415 8812 8424
rect 8760 8381 8769 8415
rect 8769 8381 8803 8415
rect 8803 8381 8812 8415
rect 8944 8415 8996 8424
rect 8760 8372 8812 8381
rect 8944 8381 8953 8415
rect 8953 8381 8987 8415
rect 8987 8381 8996 8415
rect 8944 8372 8996 8381
rect 9312 8483 9364 8492
rect 9312 8449 9321 8483
rect 9321 8449 9355 8483
rect 9355 8449 9364 8483
rect 9312 8440 9364 8449
rect 9496 8415 9548 8424
rect 5908 8236 5960 8288
rect 6552 8279 6604 8288
rect 6552 8245 6561 8279
rect 6561 8245 6595 8279
rect 6595 8245 6604 8279
rect 6552 8236 6604 8245
rect 9496 8381 9505 8415
rect 9505 8381 9539 8415
rect 9539 8381 9548 8415
rect 9496 8372 9548 8381
rect 10140 8508 10192 8560
rect 10508 8551 10560 8560
rect 9404 8304 9456 8356
rect 10048 8372 10100 8424
rect 10508 8517 10517 8551
rect 10517 8517 10551 8551
rect 10551 8517 10560 8551
rect 10508 8508 10560 8517
rect 11796 8508 11848 8560
rect 10692 8440 10744 8492
rect 10876 8372 10928 8424
rect 12808 8440 12860 8492
rect 12532 8372 12584 8424
rect 12900 8372 12952 8424
rect 10140 8347 10192 8356
rect 10140 8313 10149 8347
rect 10149 8313 10183 8347
rect 10183 8313 10192 8347
rect 10140 8304 10192 8313
rect 10232 8304 10284 8356
rect 9772 8236 9824 8288
rect 10416 8236 10468 8288
rect 12072 8279 12124 8288
rect 12072 8245 12081 8279
rect 12081 8245 12115 8279
rect 12115 8245 12124 8279
rect 12072 8236 12124 8245
rect 12624 8304 12676 8356
rect 8246 8134 8298 8186
rect 8310 8134 8362 8186
rect 8374 8134 8426 8186
rect 8438 8134 8490 8186
rect 4160 8032 4212 8084
rect 5632 8075 5684 8084
rect 5632 8041 5641 8075
rect 5641 8041 5675 8075
rect 5675 8041 5684 8075
rect 5632 8032 5684 8041
rect 6184 8075 6236 8084
rect 6184 8041 6193 8075
rect 6193 8041 6227 8075
rect 6227 8041 6236 8075
rect 6184 8032 6236 8041
rect 6644 8032 6696 8084
rect 3884 7964 3936 8016
rect 1400 7896 1452 7948
rect 2412 7896 2464 7948
rect 3332 7939 3384 7948
rect 3332 7905 3341 7939
rect 3341 7905 3375 7939
rect 3375 7905 3384 7939
rect 3332 7896 3384 7905
rect 3976 7896 4028 7948
rect 5356 7939 5408 7948
rect 5356 7905 5365 7939
rect 5365 7905 5399 7939
rect 5399 7905 5408 7939
rect 7748 7964 7800 8016
rect 9680 8032 9732 8084
rect 10140 8032 10192 8084
rect 10416 8032 10468 8084
rect 10232 7964 10284 8016
rect 10508 8007 10560 8016
rect 10508 7973 10517 8007
rect 10517 7973 10551 8007
rect 10551 7973 10560 8007
rect 10508 7964 10560 7973
rect 11796 7964 11848 8016
rect 13360 7964 13412 8016
rect 5816 7939 5868 7948
rect 5356 7896 5408 7905
rect 5816 7905 5825 7939
rect 5825 7905 5859 7939
rect 5859 7905 5868 7939
rect 5816 7896 5868 7905
rect 6920 7896 6972 7948
rect 7196 7939 7248 7948
rect 7196 7905 7205 7939
rect 7205 7905 7239 7939
rect 7239 7905 7248 7939
rect 7196 7896 7248 7905
rect 7380 7896 7432 7948
rect 8116 7896 8168 7948
rect 9128 7939 9180 7948
rect 9128 7905 9137 7939
rect 9137 7905 9171 7939
rect 9171 7905 9180 7939
rect 9128 7896 9180 7905
rect 6828 7871 6880 7880
rect 6828 7837 6837 7871
rect 6837 7837 6871 7871
rect 6871 7837 6880 7871
rect 6828 7828 6880 7837
rect 7840 7871 7892 7880
rect 7840 7837 7849 7871
rect 7849 7837 7883 7871
rect 7883 7837 7892 7871
rect 7840 7828 7892 7837
rect 2964 7803 3016 7812
rect 2964 7769 2973 7803
rect 2973 7769 3007 7803
rect 3007 7769 3016 7803
rect 2964 7760 3016 7769
rect 6368 7760 6420 7812
rect 5908 7692 5960 7744
rect 7288 7735 7340 7744
rect 7288 7701 7297 7735
rect 7297 7701 7331 7735
rect 7331 7701 7340 7735
rect 7288 7692 7340 7701
rect 8024 7692 8076 7744
rect 10048 7896 10100 7948
rect 12072 7896 12124 7948
rect 13268 7939 13320 7948
rect 13268 7905 13277 7939
rect 13277 7905 13311 7939
rect 13311 7905 13320 7939
rect 13268 7896 13320 7905
rect 10232 7871 10284 7880
rect 10232 7837 10241 7871
rect 10241 7837 10275 7871
rect 10275 7837 10284 7871
rect 10232 7828 10284 7837
rect 10600 7828 10652 7880
rect 10876 7692 10928 7744
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 12246 7590 12298 7642
rect 12310 7590 12362 7642
rect 12374 7590 12426 7642
rect 12438 7590 12490 7642
rect 5816 7488 5868 7540
rect 7656 7488 7708 7540
rect 6828 7420 6880 7472
rect 1400 7352 1452 7404
rect 2780 7352 2832 7404
rect 5264 7395 5316 7404
rect 5264 7361 5273 7395
rect 5273 7361 5307 7395
rect 5307 7361 5316 7395
rect 5264 7352 5316 7361
rect 5448 7352 5500 7404
rect 2964 7327 3016 7336
rect 2964 7293 2973 7327
rect 2973 7293 3007 7327
rect 3007 7293 3016 7327
rect 2964 7284 3016 7293
rect 3332 7284 3384 7336
rect 2504 7216 2556 7268
rect 3516 7284 3568 7336
rect 4344 7284 4396 7336
rect 3792 7216 3844 7268
rect 4528 7259 4580 7268
rect 4528 7225 4537 7259
rect 4537 7225 4571 7259
rect 4571 7225 4580 7259
rect 4528 7216 4580 7225
rect 5080 7216 5132 7268
rect 5632 7216 5684 7268
rect 1676 7191 1728 7200
rect 1676 7157 1685 7191
rect 1685 7157 1719 7191
rect 1719 7157 1728 7191
rect 1676 7148 1728 7157
rect 4620 7148 4672 7200
rect 6552 7284 6604 7336
rect 9128 7488 9180 7540
rect 8116 7420 8168 7472
rect 8208 7420 8260 7472
rect 6736 7216 6788 7268
rect 7380 7216 7432 7268
rect 7656 7216 7708 7268
rect 9036 7284 9088 7336
rect 10876 7488 10928 7540
rect 9496 7463 9548 7472
rect 9496 7429 9505 7463
rect 9505 7429 9539 7463
rect 9539 7429 9548 7463
rect 9496 7420 9548 7429
rect 13360 7420 13412 7472
rect 9956 7352 10008 7404
rect 10784 7395 10836 7404
rect 9772 7284 9824 7336
rect 10784 7361 10793 7395
rect 10793 7361 10827 7395
rect 10827 7361 10836 7395
rect 10784 7352 10836 7361
rect 12992 7352 13044 7404
rect 12072 7327 12124 7336
rect 12072 7293 12081 7327
rect 12081 7293 12115 7327
rect 12115 7293 12124 7327
rect 12072 7284 12124 7293
rect 12440 7284 12492 7336
rect 8668 7148 8720 7200
rect 8760 7148 8812 7200
rect 9864 7216 9916 7268
rect 11244 7259 11296 7268
rect 11244 7225 11253 7259
rect 11253 7225 11287 7259
rect 11287 7225 11296 7259
rect 11244 7216 11296 7225
rect 9680 7148 9732 7200
rect 9956 7191 10008 7200
rect 9956 7157 9965 7191
rect 9965 7157 9999 7191
rect 9999 7157 10008 7191
rect 9956 7148 10008 7157
rect 10048 7148 10100 7200
rect 8246 7046 8298 7098
rect 8310 7046 8362 7098
rect 8374 7046 8426 7098
rect 8438 7046 8490 7098
rect 4068 6944 4120 6996
rect 7012 6944 7064 6996
rect 7840 6944 7892 6996
rect 2504 6919 2556 6928
rect 2504 6885 2513 6919
rect 2513 6885 2547 6919
rect 2547 6885 2556 6919
rect 2504 6876 2556 6885
rect 7472 6876 7524 6928
rect 8760 6944 8812 6996
rect 1400 6808 1452 6860
rect 2136 6808 2188 6860
rect 2780 6808 2832 6860
rect 3884 6851 3936 6860
rect 3884 6817 3893 6851
rect 3893 6817 3927 6851
rect 3927 6817 3936 6851
rect 3884 6808 3936 6817
rect 4344 6851 4396 6860
rect 4344 6817 4353 6851
rect 4353 6817 4387 6851
rect 4387 6817 4396 6851
rect 4344 6808 4396 6817
rect 5632 6808 5684 6860
rect 6184 6808 6236 6860
rect 6460 6808 6512 6860
rect 11244 6919 11296 6928
rect 2044 6740 2096 6792
rect 8208 6808 8260 6860
rect 8760 6808 8812 6860
rect 11244 6885 11253 6919
rect 11253 6885 11287 6919
rect 11287 6885 11296 6919
rect 11244 6876 11296 6885
rect 12072 6876 12124 6928
rect 3516 6647 3568 6656
rect 3516 6613 3525 6647
rect 3525 6613 3559 6647
rect 3559 6613 3568 6647
rect 3516 6604 3568 6613
rect 5816 6715 5868 6724
rect 5816 6681 5825 6715
rect 5825 6681 5859 6715
rect 5859 6681 5868 6715
rect 5816 6672 5868 6681
rect 8668 6740 8720 6792
rect 9404 6740 9456 6792
rect 10784 6808 10836 6860
rect 10968 6740 11020 6792
rect 12716 6740 12768 6792
rect 13084 6783 13136 6792
rect 13084 6749 13093 6783
rect 13093 6749 13127 6783
rect 13127 6749 13136 6783
rect 13084 6740 13136 6749
rect 8484 6672 8536 6724
rect 5448 6604 5500 6656
rect 7196 6604 7248 6656
rect 7380 6604 7432 6656
rect 9128 6672 9180 6724
rect 11428 6672 11480 6724
rect 11520 6672 11572 6724
rect 9036 6604 9088 6656
rect 9496 6604 9548 6656
rect 10048 6604 10100 6656
rect 10508 6604 10560 6656
rect 11704 6604 11756 6656
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 12246 6502 12298 6554
rect 12310 6502 12362 6554
rect 12374 6502 12426 6554
rect 12438 6502 12490 6554
rect 8116 6400 8168 6452
rect 2136 6332 2188 6384
rect 2872 6332 2924 6384
rect 5816 6332 5868 6384
rect 5908 6332 5960 6384
rect 7564 6332 7616 6384
rect 7656 6332 7708 6384
rect 1400 6307 1452 6316
rect 1400 6273 1409 6307
rect 1409 6273 1443 6307
rect 1443 6273 1452 6307
rect 1400 6264 1452 6273
rect 1676 6264 1728 6316
rect 1584 6196 1636 6248
rect 3884 6264 3936 6316
rect 5264 6307 5316 6316
rect 2504 6239 2556 6248
rect 2504 6205 2513 6239
rect 2513 6205 2547 6239
rect 2547 6205 2556 6239
rect 2504 6196 2556 6205
rect 5264 6273 5273 6307
rect 5273 6273 5307 6307
rect 5307 6273 5316 6307
rect 5264 6264 5316 6273
rect 5448 6307 5500 6316
rect 5448 6273 5457 6307
rect 5457 6273 5491 6307
rect 5491 6273 5500 6307
rect 5448 6264 5500 6273
rect 7932 6332 7984 6384
rect 8208 6332 8260 6384
rect 3332 6128 3384 6180
rect 5540 6196 5592 6248
rect 7012 6196 7064 6248
rect 7196 6196 7248 6248
rect 7288 6196 7340 6248
rect 7840 6239 7892 6248
rect 7840 6205 7849 6239
rect 7849 6205 7883 6239
rect 7883 6205 7892 6239
rect 8024 6239 8076 6248
rect 7840 6196 7892 6205
rect 8024 6205 8033 6239
rect 8033 6205 8067 6239
rect 8067 6205 8076 6239
rect 8024 6196 8076 6205
rect 8668 6196 8720 6248
rect 9956 6332 10008 6384
rect 9128 6239 9180 6248
rect 9128 6205 9137 6239
rect 9137 6205 9171 6239
rect 9171 6205 9180 6239
rect 9128 6196 9180 6205
rect 9036 6128 9088 6180
rect 9864 6239 9916 6248
rect 9864 6205 9873 6239
rect 9873 6205 9907 6239
rect 9907 6205 9916 6239
rect 9864 6196 9916 6205
rect 10508 6239 10560 6248
rect 10508 6205 10517 6239
rect 10517 6205 10551 6239
rect 10551 6205 10560 6239
rect 10508 6196 10560 6205
rect 12716 6264 12768 6316
rect 13268 6264 13320 6316
rect 12900 6239 12952 6248
rect 12900 6205 12909 6239
rect 12909 6205 12943 6239
rect 12943 6205 12952 6239
rect 12900 6196 12952 6205
rect 10692 6171 10744 6180
rect 10692 6137 10701 6171
rect 10701 6137 10735 6171
rect 10735 6137 10744 6171
rect 10692 6128 10744 6137
rect 10784 6171 10836 6180
rect 10784 6137 10793 6171
rect 10793 6137 10827 6171
rect 10827 6137 10836 6171
rect 10784 6128 10836 6137
rect 7748 6060 7800 6112
rect 9864 6060 9916 6112
rect 9956 6060 10008 6112
rect 11152 6060 11204 6112
rect 12808 6060 12860 6112
rect 13176 6103 13228 6112
rect 13176 6069 13185 6103
rect 13185 6069 13219 6103
rect 13219 6069 13228 6103
rect 13176 6060 13228 6069
rect 8246 5958 8298 6010
rect 8310 5958 8362 6010
rect 8374 5958 8426 6010
rect 8438 5958 8490 6010
rect 1400 5899 1452 5908
rect 1400 5865 1409 5899
rect 1409 5865 1443 5899
rect 1443 5865 1452 5899
rect 1400 5856 1452 5865
rect 1860 5899 1912 5908
rect 1860 5865 1869 5899
rect 1869 5865 1903 5899
rect 1903 5865 1912 5899
rect 1860 5856 1912 5865
rect 3056 5788 3108 5840
rect 4804 5788 4856 5840
rect 6736 5856 6788 5908
rect 6184 5788 6236 5840
rect 6368 5788 6420 5840
rect 7196 5788 7248 5840
rect 7932 5788 7984 5840
rect 3332 5763 3384 5772
rect 3332 5729 3341 5763
rect 3341 5729 3375 5763
rect 3375 5729 3384 5763
rect 3332 5720 3384 5729
rect 3516 5720 3568 5772
rect 4712 5720 4764 5772
rect 5632 5763 5684 5772
rect 2044 5695 2096 5704
rect 2044 5661 2053 5695
rect 2053 5661 2087 5695
rect 2087 5661 2096 5695
rect 2044 5652 2096 5661
rect 2872 5695 2924 5704
rect 2872 5661 2881 5695
rect 2881 5661 2915 5695
rect 2915 5661 2924 5695
rect 2872 5652 2924 5661
rect 5632 5729 5641 5763
rect 5641 5729 5675 5763
rect 5675 5729 5684 5763
rect 5632 5720 5684 5729
rect 7840 5652 7892 5704
rect 9036 5788 9088 5840
rect 8760 5720 8812 5772
rect 10784 5856 10836 5908
rect 10968 5899 11020 5908
rect 10968 5865 10977 5899
rect 10977 5865 11011 5899
rect 11011 5865 11020 5899
rect 10968 5856 11020 5865
rect 9772 5788 9824 5840
rect 9864 5763 9916 5772
rect 8668 5652 8720 5704
rect 9864 5729 9873 5763
rect 9873 5729 9907 5763
rect 9907 5729 9916 5763
rect 9864 5720 9916 5729
rect 10692 5788 10744 5840
rect 11244 5788 11296 5840
rect 11704 5831 11756 5840
rect 11704 5797 11713 5831
rect 11713 5797 11747 5831
rect 11747 5797 11756 5831
rect 11704 5788 11756 5797
rect 13176 5788 13228 5840
rect 9772 5652 9824 5704
rect 5540 5516 5592 5568
rect 7380 5559 7432 5568
rect 7380 5525 7389 5559
rect 7389 5525 7423 5559
rect 7423 5525 7432 5559
rect 7380 5516 7432 5525
rect 8024 5559 8076 5568
rect 8024 5525 8033 5559
rect 8033 5525 8067 5559
rect 8067 5525 8076 5559
rect 8024 5516 8076 5525
rect 8484 5559 8536 5568
rect 8484 5525 8493 5559
rect 8493 5525 8527 5559
rect 8527 5525 8536 5559
rect 8484 5516 8536 5525
rect 9036 5584 9088 5636
rect 9864 5584 9916 5636
rect 9588 5516 9640 5568
rect 10232 5652 10284 5704
rect 11520 5516 11572 5568
rect 13176 5559 13228 5568
rect 13176 5525 13185 5559
rect 13185 5525 13219 5559
rect 13219 5525 13228 5559
rect 13176 5516 13228 5525
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 12246 5414 12298 5466
rect 12310 5414 12362 5466
rect 12374 5414 12426 5466
rect 12438 5414 12490 5466
rect 5632 5312 5684 5364
rect 6000 5312 6052 5364
rect 7472 5312 7524 5364
rect 8760 5355 8812 5364
rect 4344 5176 4396 5228
rect 1584 5151 1636 5160
rect 1584 5117 1593 5151
rect 1593 5117 1627 5151
rect 1627 5117 1636 5151
rect 1584 5108 1636 5117
rect 4068 5108 4120 5160
rect 4620 5108 4672 5160
rect 6000 5151 6052 5160
rect 6000 5117 6009 5151
rect 6009 5117 6043 5151
rect 6043 5117 6052 5151
rect 8024 5176 8076 5228
rect 8760 5321 8769 5355
rect 8769 5321 8803 5355
rect 8803 5321 8812 5355
rect 8760 5312 8812 5321
rect 9404 5176 9456 5228
rect 10232 5312 10284 5364
rect 10784 5312 10836 5364
rect 9772 5219 9824 5228
rect 9772 5185 9781 5219
rect 9781 5185 9815 5219
rect 9815 5185 9824 5219
rect 9772 5176 9824 5185
rect 12440 5176 12492 5228
rect 13176 5219 13228 5228
rect 13176 5185 13185 5219
rect 13185 5185 13219 5219
rect 13219 5185 13228 5219
rect 13176 5176 13228 5185
rect 6000 5108 6052 5117
rect 11888 5151 11940 5160
rect 11888 5117 11897 5151
rect 11897 5117 11931 5151
rect 11931 5117 11940 5151
rect 11888 5108 11940 5117
rect 3608 5083 3660 5092
rect 3608 5049 3617 5083
rect 3617 5049 3651 5083
rect 3651 5049 3660 5083
rect 3608 5040 3660 5049
rect 5724 5083 5776 5092
rect 5724 5049 5733 5083
rect 5733 5049 5767 5083
rect 5767 5049 5776 5083
rect 5724 5040 5776 5049
rect 5816 5040 5868 5092
rect 11152 5040 11204 5092
rect 13084 5083 13136 5092
rect 13084 5049 13093 5083
rect 13093 5049 13127 5083
rect 13127 5049 13136 5083
rect 13084 5040 13136 5049
rect 2136 5015 2188 5024
rect 2136 4981 2145 5015
rect 2145 4981 2179 5015
rect 2179 4981 2188 5015
rect 2136 4972 2188 4981
rect 6368 4972 6420 5024
rect 6552 5015 6604 5024
rect 6552 4981 6561 5015
rect 6561 4981 6595 5015
rect 6595 4981 6604 5015
rect 6552 4972 6604 4981
rect 11796 5015 11848 5024
rect 11796 4981 11805 5015
rect 11805 4981 11839 5015
rect 11839 4981 11848 5015
rect 11796 4972 11848 4981
rect 8246 4870 8298 4922
rect 8310 4870 8362 4922
rect 8374 4870 8426 4922
rect 8438 4870 8490 4922
rect 2044 4675 2096 4684
rect 2044 4641 2053 4675
rect 2053 4641 2087 4675
rect 2087 4641 2096 4675
rect 2044 4632 2096 4641
rect 2136 4632 2188 4684
rect 3608 4768 3660 4820
rect 4160 4768 4212 4820
rect 1952 4564 2004 4616
rect 2964 4607 3016 4616
rect 2964 4573 2973 4607
rect 2973 4573 3007 4607
rect 3007 4573 3016 4607
rect 2964 4564 3016 4573
rect 3424 4632 3476 4684
rect 5724 4768 5776 4820
rect 5356 4700 5408 4752
rect 4160 4675 4212 4684
rect 4160 4641 4164 4675
rect 4164 4641 4198 4675
rect 4198 4641 4212 4675
rect 4344 4675 4396 4684
rect 4160 4632 4212 4641
rect 4344 4641 4353 4675
rect 4353 4641 4387 4675
rect 4387 4641 4396 4675
rect 4344 4632 4396 4641
rect 6736 4700 6788 4752
rect 3884 4564 3936 4616
rect 2872 4428 2924 4480
rect 4620 4496 4672 4548
rect 4896 4564 4948 4616
rect 5724 4564 5776 4616
rect 6368 4675 6420 4684
rect 6368 4641 6377 4675
rect 6377 4641 6411 4675
rect 6411 4641 6420 4675
rect 6368 4632 6420 4641
rect 6828 4675 6880 4684
rect 6828 4641 6837 4675
rect 6837 4641 6871 4675
rect 6871 4641 6880 4675
rect 6828 4632 6880 4641
rect 7380 4632 7432 4684
rect 7656 4632 7708 4684
rect 8852 4768 8904 4820
rect 13084 4768 13136 4820
rect 9128 4743 9180 4752
rect 9128 4709 9137 4743
rect 9137 4709 9171 4743
rect 9171 4709 9180 4743
rect 9128 4700 9180 4709
rect 12808 4700 12860 4752
rect 8668 4632 8720 4684
rect 8852 4632 8904 4684
rect 9864 4675 9916 4684
rect 7012 4564 7064 4616
rect 5540 4496 5592 4548
rect 7380 4471 7432 4480
rect 7380 4437 7389 4471
rect 7389 4437 7423 4471
rect 7423 4437 7432 4471
rect 7380 4428 7432 4437
rect 8116 4428 8168 4480
rect 8392 4428 8444 4480
rect 8760 4564 8812 4616
rect 9496 4607 9548 4616
rect 9496 4573 9505 4607
rect 9505 4573 9539 4607
rect 9539 4573 9548 4607
rect 9496 4564 9548 4573
rect 9864 4641 9873 4675
rect 9873 4641 9907 4675
rect 9907 4641 9916 4675
rect 9864 4632 9916 4641
rect 10600 4632 10652 4684
rect 11060 4632 11112 4684
rect 11520 4675 11572 4684
rect 11520 4641 11529 4675
rect 11529 4641 11563 4675
rect 11563 4641 11572 4675
rect 11520 4632 11572 4641
rect 10140 4607 10192 4616
rect 10140 4573 10149 4607
rect 10149 4573 10183 4607
rect 10183 4573 10192 4607
rect 10140 4564 10192 4573
rect 10692 4607 10744 4616
rect 10692 4573 10701 4607
rect 10701 4573 10735 4607
rect 10735 4573 10744 4607
rect 10692 4564 10744 4573
rect 12440 4564 12492 4616
rect 9772 4496 9824 4548
rect 10048 4496 10100 4548
rect 8760 4428 8812 4480
rect 11060 4471 11112 4480
rect 11060 4437 11069 4471
rect 11069 4437 11103 4471
rect 11103 4437 11112 4471
rect 11060 4428 11112 4437
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 12246 4326 12298 4378
rect 12310 4326 12362 4378
rect 12374 4326 12426 4378
rect 12438 4326 12490 4378
rect 2872 4224 2924 4276
rect 2044 4156 2096 4208
rect 4436 4156 4488 4208
rect 11888 4156 11940 4208
rect 480 4088 532 4140
rect 1492 4088 1544 4140
rect 8116 4131 8168 4140
rect 1768 4063 1820 4072
rect 1768 4029 1777 4063
rect 1777 4029 1811 4063
rect 1811 4029 1820 4063
rect 1768 4020 1820 4029
rect 1952 4063 2004 4072
rect 1952 4029 1961 4063
rect 1961 4029 1995 4063
rect 1995 4029 2004 4063
rect 1952 4020 2004 4029
rect 2136 4063 2188 4072
rect 2136 4029 2146 4063
rect 2146 4029 2180 4063
rect 2180 4029 2188 4063
rect 2964 4063 3016 4072
rect 2136 4020 2188 4029
rect 2964 4029 2973 4063
rect 2973 4029 3007 4063
rect 3007 4029 3016 4063
rect 2964 4020 3016 4029
rect 3884 4020 3936 4072
rect 6000 4020 6052 4072
rect 6736 4063 6788 4072
rect 6736 4029 6740 4063
rect 6740 4029 6774 4063
rect 6774 4029 6788 4063
rect 6736 4020 6788 4029
rect 7104 4063 7156 4072
rect 7104 4029 7113 4063
rect 7113 4029 7147 4063
rect 7147 4029 7156 4063
rect 7104 4020 7156 4029
rect 7380 4020 7432 4072
rect 8116 4097 8125 4131
rect 8125 4097 8159 4131
rect 8159 4097 8168 4131
rect 8116 4088 8168 4097
rect 8760 4088 8812 4140
rect 9772 4088 9824 4140
rect 11244 4131 11296 4140
rect 11244 4097 11253 4131
rect 11253 4097 11287 4131
rect 11287 4097 11296 4131
rect 11244 4088 11296 4097
rect 8392 4020 8444 4072
rect 8576 4020 8628 4072
rect 9404 4020 9456 4072
rect 11796 4020 11848 4072
rect 12900 4156 12952 4208
rect 12900 4020 12952 4072
rect 13084 4020 13136 4072
rect 3332 3952 3384 4004
rect 5632 3995 5684 4004
rect 2228 3884 2280 3936
rect 3424 3927 3476 3936
rect 3424 3893 3433 3927
rect 3433 3893 3467 3927
rect 3467 3893 3476 3927
rect 3424 3884 3476 3893
rect 3884 3884 3936 3936
rect 5632 3961 5641 3995
rect 5641 3961 5675 3995
rect 5675 3961 5684 3995
rect 5632 3952 5684 3961
rect 6368 3952 6420 4004
rect 6828 3995 6880 4004
rect 6828 3961 6837 3995
rect 6837 3961 6871 3995
rect 6871 3961 6880 3995
rect 6828 3952 6880 3961
rect 7012 3952 7064 4004
rect 8760 3995 8812 4004
rect 8760 3961 8769 3995
rect 8769 3961 8803 3995
rect 8803 3961 8812 3995
rect 8760 3952 8812 3961
rect 12072 3995 12124 4004
rect 4620 3884 4672 3936
rect 4712 3884 4764 3936
rect 4988 3884 5040 3936
rect 6276 3884 6328 3936
rect 6736 3884 6788 3936
rect 12072 3961 12081 3995
rect 12081 3961 12115 3995
rect 12115 3961 12124 3995
rect 12072 3952 12124 3961
rect 12716 3927 12768 3936
rect 12716 3893 12725 3927
rect 12725 3893 12759 3927
rect 12759 3893 12768 3927
rect 12716 3884 12768 3893
rect 8246 3782 8298 3834
rect 8310 3782 8362 3834
rect 8374 3782 8426 3834
rect 8438 3782 8490 3834
rect 5356 3723 5408 3732
rect 5356 3689 5365 3723
rect 5365 3689 5399 3723
rect 5399 3689 5408 3723
rect 5356 3680 5408 3689
rect 5448 3723 5500 3732
rect 5448 3689 5457 3723
rect 5457 3689 5491 3723
rect 5491 3689 5500 3723
rect 5632 3723 5684 3732
rect 5448 3680 5500 3689
rect 5632 3689 5641 3723
rect 5641 3689 5675 3723
rect 5675 3689 5684 3723
rect 5632 3680 5684 3689
rect 1492 3587 1544 3596
rect 1492 3553 1501 3587
rect 1501 3553 1535 3587
rect 1535 3553 1544 3587
rect 1492 3544 1544 3553
rect 1676 3587 1728 3596
rect 1676 3553 1685 3587
rect 1685 3553 1719 3587
rect 1719 3553 1728 3587
rect 1676 3544 1728 3553
rect 1860 3544 1912 3596
rect 2044 3544 2096 3596
rect 2228 3587 2280 3596
rect 2228 3553 2237 3587
rect 2237 3553 2271 3587
rect 2271 3553 2280 3587
rect 2228 3544 2280 3553
rect 4620 3612 4672 3664
rect 9128 3680 9180 3732
rect 3056 3544 3108 3596
rect 4528 3587 4580 3596
rect 4528 3553 4537 3587
rect 4537 3553 4571 3587
rect 4571 3553 4580 3587
rect 4528 3544 4580 3553
rect 1768 3408 1820 3460
rect 3332 3476 3384 3528
rect 4436 3476 4488 3528
rect 5540 3587 5592 3596
rect 5540 3553 5549 3587
rect 5549 3553 5583 3587
rect 5583 3553 5592 3587
rect 5540 3544 5592 3553
rect 5908 3544 5960 3596
rect 6552 3544 6604 3596
rect 7012 3612 7064 3664
rect 7104 3587 7156 3596
rect 7104 3553 7113 3587
rect 7113 3553 7147 3587
rect 7147 3553 7156 3587
rect 7104 3544 7156 3553
rect 7472 3587 7524 3596
rect 7472 3553 7481 3587
rect 7481 3553 7515 3587
rect 7515 3553 7524 3587
rect 7472 3544 7524 3553
rect 7564 3544 7616 3596
rect 8300 3612 8352 3664
rect 8392 3587 8444 3596
rect 8392 3553 8401 3587
rect 8401 3553 8435 3587
rect 8435 3553 8444 3587
rect 8392 3544 8444 3553
rect 8576 3587 8628 3596
rect 8576 3553 8585 3587
rect 8585 3553 8619 3587
rect 8619 3553 8628 3587
rect 8576 3544 8628 3553
rect 10140 3680 10192 3732
rect 11060 3680 11112 3732
rect 10600 3587 10652 3596
rect 5632 3476 5684 3528
rect 7656 3476 7708 3528
rect 5816 3408 5868 3460
rect 8760 3476 8812 3528
rect 9496 3476 9548 3528
rect 5448 3340 5500 3392
rect 8392 3408 8444 3460
rect 8944 3340 8996 3392
rect 9312 3340 9364 3392
rect 10600 3553 10609 3587
rect 10609 3553 10643 3587
rect 10643 3553 10652 3587
rect 10600 3544 10652 3553
rect 10692 3544 10744 3596
rect 10968 3587 11020 3596
rect 10968 3553 10978 3587
rect 10978 3553 11012 3587
rect 11012 3553 11020 3587
rect 11152 3587 11204 3596
rect 10968 3544 11020 3553
rect 11152 3553 11161 3587
rect 11161 3553 11195 3587
rect 11195 3553 11204 3587
rect 11152 3544 11204 3553
rect 12716 3680 12768 3732
rect 12808 3612 12860 3664
rect 11520 3519 11572 3528
rect 11520 3485 11529 3519
rect 11529 3485 11563 3519
rect 11563 3485 11572 3519
rect 11796 3519 11848 3528
rect 11520 3476 11572 3485
rect 11796 3485 11805 3519
rect 11805 3485 11839 3519
rect 11839 3485 11848 3519
rect 11796 3476 11848 3485
rect 12164 3476 12216 3528
rect 12900 3340 12952 3392
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 12246 3238 12298 3290
rect 12310 3238 12362 3290
rect 12374 3238 12426 3290
rect 12438 3238 12490 3290
rect 4620 3136 4672 3188
rect 6552 3136 6604 3188
rect 7472 3136 7524 3188
rect 7564 3179 7616 3188
rect 7564 3145 7573 3179
rect 7573 3145 7607 3179
rect 7607 3145 7616 3179
rect 7564 3136 7616 3145
rect 8392 3136 8444 3188
rect 1952 3111 2004 3120
rect 1952 3077 1961 3111
rect 1961 3077 1995 3111
rect 1995 3077 2004 3111
rect 1952 3068 2004 3077
rect 5540 3111 5592 3120
rect 1584 3000 1636 3052
rect 4068 3043 4120 3052
rect 1400 2932 1452 2984
rect 1676 2932 1728 2984
rect 4068 3009 4077 3043
rect 4077 3009 4111 3043
rect 4111 3009 4120 3043
rect 4068 3000 4120 3009
rect 5540 3077 5549 3111
rect 5549 3077 5583 3111
rect 5583 3077 5592 3111
rect 5540 3068 5592 3077
rect 5632 3068 5684 3120
rect 9312 3111 9364 3120
rect 1492 2864 1544 2916
rect 1952 2864 2004 2916
rect 3792 2907 3844 2916
rect 3792 2873 3801 2907
rect 3801 2873 3835 2907
rect 3835 2873 3844 2907
rect 3792 2864 3844 2873
rect 2504 2796 2556 2848
rect 3424 2796 3476 2848
rect 4712 2932 4764 2984
rect 5908 2975 5960 2984
rect 4804 2839 4856 2848
rect 4804 2805 4813 2839
rect 4813 2805 4847 2839
rect 4847 2805 4856 2839
rect 4804 2796 4856 2805
rect 5908 2941 5917 2975
rect 5917 2941 5951 2975
rect 5951 2941 5960 2975
rect 5908 2932 5960 2941
rect 6276 2932 6328 2984
rect 6736 2975 6788 2984
rect 6736 2941 6745 2975
rect 6745 2941 6779 2975
rect 6779 2941 6788 2975
rect 6736 2932 6788 2941
rect 7656 2932 7708 2984
rect 9312 3077 9321 3111
rect 9321 3077 9355 3111
rect 9355 3077 9364 3111
rect 9312 3068 9364 3077
rect 9864 3136 9916 3188
rect 11060 3136 11112 3188
rect 11796 3179 11848 3188
rect 11796 3145 11805 3179
rect 11805 3145 11839 3179
rect 11839 3145 11848 3179
rect 11796 3136 11848 3145
rect 12808 3136 12860 3188
rect 12992 3136 13044 3188
rect 12532 3068 12584 3120
rect 9404 3043 9456 3052
rect 9404 3009 9413 3043
rect 9413 3009 9447 3043
rect 9447 3009 9456 3043
rect 9404 3000 9456 3009
rect 8852 2975 8904 2984
rect 8852 2941 8861 2975
rect 8861 2941 8895 2975
rect 8895 2941 8904 2975
rect 8852 2932 8904 2941
rect 8944 2932 8996 2984
rect 9128 2932 9180 2984
rect 9956 2975 10008 2984
rect 9956 2941 9960 2975
rect 9960 2941 9994 2975
rect 9994 2941 10008 2975
rect 9956 2932 10008 2941
rect 10324 2975 10376 2984
rect 10324 2941 10333 2975
rect 10333 2941 10367 2975
rect 10367 2941 10376 2975
rect 10324 2932 10376 2941
rect 11244 3000 11296 3052
rect 11704 3000 11756 3052
rect 11888 2975 11940 2984
rect 11888 2941 11937 2975
rect 11937 2941 11940 2975
rect 11888 2932 11940 2941
rect 12808 2975 12860 2984
rect 12808 2941 12817 2975
rect 12817 2941 12851 2975
rect 12851 2941 12860 2975
rect 12808 2932 12860 2941
rect 13084 2932 13136 2984
rect 13268 2975 13320 2984
rect 13268 2941 13277 2975
rect 13277 2941 13311 2975
rect 13311 2941 13320 2975
rect 13268 2932 13320 2941
rect 8576 2907 8628 2916
rect 8576 2873 8585 2907
rect 8585 2873 8619 2907
rect 8619 2873 8628 2907
rect 8576 2864 8628 2873
rect 12072 2907 12124 2916
rect 5816 2796 5868 2848
rect 12072 2873 12081 2907
rect 12081 2873 12115 2907
rect 12115 2873 12124 2907
rect 12072 2864 12124 2873
rect 10232 2796 10284 2848
rect 11244 2796 11296 2848
rect 12256 2796 12308 2848
rect 8246 2694 8298 2746
rect 8310 2694 8362 2746
rect 8374 2694 8426 2746
rect 8438 2694 8490 2746
rect 4620 2592 4672 2644
rect 5356 2635 5408 2644
rect 5356 2601 5365 2635
rect 5365 2601 5399 2635
rect 5399 2601 5408 2635
rect 5356 2592 5408 2601
rect 5632 2592 5684 2644
rect 3056 2567 3108 2576
rect 3056 2533 3065 2567
rect 3065 2533 3099 2567
rect 3099 2533 3108 2567
rect 3056 2524 3108 2533
rect 1952 2456 2004 2508
rect 2320 2499 2372 2508
rect 2320 2465 2329 2499
rect 2329 2465 2363 2499
rect 2363 2465 2372 2499
rect 2320 2456 2372 2465
rect 2504 2499 2556 2508
rect 2504 2465 2513 2499
rect 2513 2465 2547 2499
rect 2547 2465 2556 2499
rect 4804 2524 4856 2576
rect 6368 2592 6420 2644
rect 7656 2592 7708 2644
rect 6276 2524 6328 2576
rect 2504 2456 2556 2465
rect 3332 2456 3384 2508
rect 4160 2499 4212 2508
rect 4160 2465 4164 2499
rect 4164 2465 4198 2499
rect 4198 2465 4212 2499
rect 4160 2456 4212 2465
rect 5172 2499 5224 2508
rect 5172 2465 5181 2499
rect 5181 2465 5215 2499
rect 5215 2465 5224 2499
rect 5172 2456 5224 2465
rect 5356 2456 5408 2508
rect 5632 2456 5684 2508
rect 6184 2499 6236 2508
rect 6184 2465 6193 2499
rect 6193 2465 6227 2499
rect 6227 2465 6236 2499
rect 6184 2456 6236 2465
rect 2320 2320 2372 2372
rect 3332 2320 3384 2372
rect 3792 2320 3844 2372
rect 4160 2320 4212 2372
rect 4620 2320 4672 2372
rect 6552 2456 6604 2508
rect 6736 2499 6788 2508
rect 6736 2465 6745 2499
rect 6745 2465 6779 2499
rect 6779 2465 6788 2499
rect 6736 2456 6788 2465
rect 8116 2499 8168 2508
rect 5724 2320 5776 2372
rect 5816 2320 5868 2372
rect 6644 2320 6696 2372
rect 8116 2465 8125 2499
rect 8125 2465 8159 2499
rect 8159 2465 8168 2499
rect 8116 2456 8168 2465
rect 8944 2524 8996 2576
rect 10692 2592 10744 2644
rect 12256 2592 12308 2644
rect 8852 2456 8904 2508
rect 9220 2456 9272 2508
rect 10324 2456 10376 2508
rect 11152 2524 11204 2576
rect 10692 2456 10744 2508
rect 11520 2524 11572 2576
rect 12624 2524 12676 2576
rect 8760 2388 8812 2440
rect 5356 2252 5408 2304
rect 5540 2252 5592 2304
rect 7564 2295 7616 2304
rect 7564 2261 7573 2295
rect 7573 2261 7607 2295
rect 7607 2261 7616 2295
rect 7564 2252 7616 2261
rect 9404 2388 9456 2440
rect 11612 2431 11664 2440
rect 11612 2397 11621 2431
rect 11621 2397 11655 2431
rect 11655 2397 11664 2431
rect 11612 2388 11664 2397
rect 11060 2320 11112 2372
rect 11796 2252 11848 2304
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 12246 2150 12298 2202
rect 12310 2150 12362 2202
rect 12374 2150 12426 2202
rect 12438 2150 12490 2202
rect 2320 2048 2372 2100
rect 4620 2048 4672 2100
rect 4252 1980 4304 2032
rect 5448 1980 5500 2032
rect 4068 1912 4120 1964
rect 4160 1912 4212 1964
rect 4804 1955 4856 1964
rect 4804 1921 4813 1955
rect 4813 1921 4847 1955
rect 4847 1921 4856 1955
rect 4804 1912 4856 1921
rect 4620 1844 4672 1896
rect 2872 1776 2924 1828
rect 5356 1844 5408 1896
rect 5632 1887 5684 1896
rect 5632 1853 5641 1887
rect 5641 1853 5675 1887
rect 5675 1853 5684 1887
rect 5632 1844 5684 1853
rect 6276 2048 6328 2100
rect 9220 2091 9272 2100
rect 5816 1912 5868 1964
rect 3976 1708 4028 1760
rect 5172 1776 5224 1828
rect 6000 1844 6052 1896
rect 6552 1844 6604 1896
rect 9220 2057 9229 2091
rect 9229 2057 9263 2091
rect 9263 2057 9272 2091
rect 9220 2048 9272 2057
rect 10324 2048 10376 2100
rect 11612 2048 11664 2100
rect 12716 2048 12768 2100
rect 8116 1912 8168 1964
rect 8576 1955 8628 1964
rect 8576 1921 8585 1955
rect 8585 1921 8619 1955
rect 8619 1921 8628 1955
rect 8576 1912 8628 1921
rect 8944 1844 8996 1896
rect 10048 1980 10100 2032
rect 11060 1980 11112 2032
rect 11888 1980 11940 2032
rect 12256 2023 12308 2032
rect 10232 1844 10284 1896
rect 10968 1819 11020 1828
rect 4620 1708 4672 1760
rect 6184 1708 6236 1760
rect 6828 1708 6880 1760
rect 9772 1708 9824 1760
rect 10048 1751 10100 1760
rect 10048 1717 10057 1751
rect 10057 1717 10091 1751
rect 10091 1717 10100 1751
rect 10048 1708 10100 1717
rect 10968 1785 10977 1819
rect 10977 1785 11011 1819
rect 11011 1785 11020 1819
rect 10968 1776 11020 1785
rect 11336 1844 11388 1896
rect 12256 1989 12265 2023
rect 12265 1989 12299 2023
rect 12299 1989 12308 2023
rect 12256 1980 12308 1989
rect 12808 1887 12860 1896
rect 12808 1853 12817 1887
rect 12817 1853 12851 1887
rect 12851 1853 12860 1887
rect 12808 1844 12860 1853
rect 12900 1844 12952 1896
rect 8246 1606 8298 1658
rect 8310 1606 8362 1658
rect 8374 1606 8426 1658
rect 8438 1606 8490 1658
rect 2872 1547 2924 1556
rect 2872 1513 2881 1547
rect 2881 1513 2915 1547
rect 2915 1513 2924 1547
rect 2872 1504 2924 1513
rect 6644 1547 6696 1556
rect 6644 1513 6653 1547
rect 6653 1513 6687 1547
rect 6687 1513 6696 1547
rect 6644 1504 6696 1513
rect 6736 1504 6788 1556
rect 8760 1547 8812 1556
rect 8760 1513 8769 1547
rect 8769 1513 8803 1547
rect 8803 1513 8812 1547
rect 8760 1504 8812 1513
rect 9772 1547 9824 1556
rect 1952 1368 2004 1420
rect 2688 1411 2740 1420
rect 2688 1377 2697 1411
rect 2697 1377 2731 1411
rect 2731 1377 2740 1411
rect 2688 1368 2740 1377
rect 3332 1411 3384 1420
rect 3332 1377 3341 1411
rect 3341 1377 3375 1411
rect 3375 1377 3384 1411
rect 3332 1368 3384 1377
rect 3976 1411 4028 1420
rect 3976 1377 3985 1411
rect 3985 1377 4019 1411
rect 4019 1377 4028 1411
rect 3976 1368 4028 1377
rect 4252 1368 4304 1420
rect 7564 1436 7616 1488
rect 9772 1513 9781 1547
rect 9781 1513 9815 1547
rect 9815 1513 9824 1547
rect 9772 1504 9824 1513
rect 12624 1504 12676 1556
rect 9404 1411 9456 1420
rect 9404 1377 9413 1411
rect 9413 1377 9447 1411
rect 9447 1377 9456 1411
rect 9404 1368 9456 1377
rect 11520 1411 11572 1420
rect 11520 1377 11529 1411
rect 11529 1377 11563 1411
rect 11563 1377 11572 1411
rect 11520 1368 11572 1377
rect 12808 1368 12860 1420
rect 4620 1343 4672 1352
rect 4160 1232 4212 1284
rect 4068 1164 4120 1216
rect 4620 1309 4629 1343
rect 4629 1309 4663 1343
rect 4663 1309 4672 1343
rect 4620 1300 4672 1309
rect 6828 1300 6880 1352
rect 12256 1300 12308 1352
rect 6184 1164 6236 1216
rect 4246 1062 4298 1114
rect 4310 1062 4362 1114
rect 4374 1062 4426 1114
rect 4438 1062 4490 1114
rect 12246 1062 12298 1114
rect 12310 1062 12362 1114
rect 12374 1062 12426 1114
rect 12438 1062 12490 1114
<< metal2 >>
rect 478 16200 534 17000
rect 1858 16200 1914 17000
rect 3238 16200 3294 17000
rect 4618 16200 4674 17000
rect 5998 16200 6054 17000
rect 6918 16200 6974 17000
rect 8298 16200 8354 17000
rect 9678 16200 9734 17000
rect 11058 16200 11114 17000
rect 12438 16200 12494 17000
rect 13818 16200 13874 17000
rect 492 11762 520 16200
rect 1872 14618 1900 16200
rect 1860 14612 1912 14618
rect 1860 14554 1912 14560
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 2044 14408 2096 14414
rect 2044 14350 2096 14356
rect 1768 14272 1820 14278
rect 1768 14214 1820 14220
rect 1780 13870 1808 14214
rect 1768 13864 1820 13870
rect 1768 13806 1820 13812
rect 1780 13394 1808 13806
rect 1768 13388 1820 13394
rect 1768 13330 1820 13336
rect 2056 12918 2084 14350
rect 2780 14340 2832 14346
rect 2780 14282 2832 14288
rect 2792 13802 2820 14282
rect 2504 13796 2556 13802
rect 2504 13738 2556 13744
rect 2780 13796 2832 13802
rect 2780 13738 2832 13744
rect 2516 13462 2544 13738
rect 2504 13456 2556 13462
rect 2504 13398 2556 13404
rect 2792 13326 2820 13738
rect 3068 13530 3096 14418
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 3056 13524 3108 13530
rect 3056 13466 3108 13472
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 2044 12912 2096 12918
rect 2044 12854 2096 12860
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1688 12345 1716 12582
rect 1674 12336 1730 12345
rect 1674 12271 1730 12280
rect 2056 12238 2084 12854
rect 2136 12640 2188 12646
rect 2136 12582 2188 12588
rect 2148 12306 2176 12582
rect 2792 12306 2820 13262
rect 2136 12300 2188 12306
rect 2136 12242 2188 12248
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 2044 12232 2096 12238
rect 2044 12174 2096 12180
rect 480 11756 532 11762
rect 480 11698 532 11704
rect 2056 11694 2084 12174
rect 2884 11778 2912 13466
rect 3056 13388 3108 13394
rect 3056 13330 3108 13336
rect 2964 13184 3016 13190
rect 2964 13126 3016 13132
rect 2976 12850 3004 13126
rect 3068 12918 3096 13330
rect 3252 12918 3280 16200
rect 4632 15706 4660 16200
rect 4620 15700 4672 15706
rect 4620 15642 4672 15648
rect 4988 15632 5040 15638
rect 4988 15574 5040 15580
rect 4896 15564 4948 15570
rect 4896 15506 4948 15512
rect 4804 15496 4856 15502
rect 4804 15438 4856 15444
rect 4068 15360 4120 15366
rect 4068 15302 4120 15308
rect 4620 15360 4672 15366
rect 4620 15302 4672 15308
rect 4080 14550 4108 15302
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 4632 14958 4660 15302
rect 4620 14952 4672 14958
rect 4620 14894 4672 14900
rect 4068 14544 4120 14550
rect 4068 14486 4120 14492
rect 4632 14482 4660 14894
rect 4816 14822 4844 15438
rect 4908 14958 4936 15506
rect 4896 14952 4948 14958
rect 4896 14894 4948 14900
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 4816 14550 4844 14758
rect 4804 14544 4856 14550
rect 4804 14486 4856 14492
rect 4620 14476 4672 14482
rect 4620 14418 4672 14424
rect 3332 14408 3384 14414
rect 3332 14350 3384 14356
rect 4066 14376 4122 14385
rect 3344 13870 3372 14350
rect 3884 14340 3936 14346
rect 4066 14311 4122 14320
rect 3884 14282 3936 14288
rect 3896 13938 3924 14282
rect 4080 14006 4108 14311
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 4068 14000 4120 14006
rect 4068 13942 4120 13948
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 3332 13864 3384 13870
rect 3332 13806 3384 13812
rect 3056 12912 3108 12918
rect 3056 12854 3108 12860
rect 3240 12912 3292 12918
rect 3240 12854 3292 12860
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 3068 12374 3096 12854
rect 3148 12776 3200 12782
rect 3148 12718 3200 12724
rect 3056 12368 3108 12374
rect 3056 12310 3108 12316
rect 3160 12170 3188 12718
rect 3148 12164 3200 12170
rect 3148 12106 3200 12112
rect 2700 11750 2912 11778
rect 2044 11688 2096 11694
rect 2044 11630 2096 11636
rect 1768 11552 1820 11558
rect 1768 11494 1820 11500
rect 1780 11218 1808 11494
rect 1768 11212 1820 11218
rect 1768 11154 1820 11160
rect 1860 10600 1912 10606
rect 1860 10542 1912 10548
rect 1872 10130 1900 10542
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1860 10124 1912 10130
rect 1860 10066 1912 10072
rect 1412 9722 1440 10066
rect 1400 9716 1452 9722
rect 1400 9658 1452 9664
rect 2056 9586 2084 11630
rect 2700 11218 2728 11750
rect 3160 11694 3188 12106
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3148 11688 3200 11694
rect 3148 11630 3200 11636
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 2780 11620 2832 11626
rect 2780 11562 2832 11568
rect 3332 11620 3384 11626
rect 3332 11562 3384 11568
rect 2412 11212 2464 11218
rect 2412 11154 2464 11160
rect 2688 11212 2740 11218
rect 2688 11154 2740 11160
rect 2424 11082 2452 11154
rect 2412 11076 2464 11082
rect 2412 11018 2464 11024
rect 2424 10674 2452 11018
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 2700 10606 2728 11154
rect 2792 10606 2820 11562
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2976 10810 3004 11086
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 2688 10600 2740 10606
rect 2688 10542 2740 10548
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2700 10130 2728 10542
rect 2964 10532 3016 10538
rect 2964 10474 3016 10480
rect 2976 10198 3004 10474
rect 2964 10192 3016 10198
rect 2964 10134 3016 10140
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 3344 10112 3372 11562
rect 3436 11354 3464 11630
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3804 11286 3832 12038
rect 3792 11280 3844 11286
rect 3792 11222 3844 11228
rect 3424 10124 3476 10130
rect 3344 10084 3424 10112
rect 3344 9722 3372 10084
rect 3424 10066 3476 10072
rect 3332 9716 3384 9722
rect 3332 9658 3384 9664
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 1492 9376 1544 9382
rect 1492 9318 1544 9324
rect 1400 8288 1452 8294
rect 1400 8230 1452 8236
rect 1412 7954 1440 8230
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 1412 7410 1440 7890
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1400 6860 1452 6866
rect 1400 6802 1452 6808
rect 1412 6322 1440 6802
rect 1400 6316 1452 6322
rect 1400 6258 1452 6264
rect 1412 5914 1440 6258
rect 1400 5908 1452 5914
rect 1400 5850 1452 5856
rect 1504 4146 1532 9318
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1780 8430 1808 8774
rect 2056 8498 2084 9522
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2136 9036 2188 9042
rect 2136 8978 2188 8984
rect 2320 9036 2372 9042
rect 2372 8996 2452 9024
rect 2320 8978 2372 8984
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 1768 8424 1820 8430
rect 1768 8366 1820 8372
rect 1860 8356 1912 8362
rect 1860 8298 1912 8304
rect 1872 8265 1900 8298
rect 1858 8256 1914 8265
rect 1858 8191 1914 8200
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 1688 6322 1716 7142
rect 2056 6798 2084 8434
rect 2148 6866 2176 8978
rect 2424 8362 2452 8996
rect 2412 8356 2464 8362
rect 2412 8298 2464 8304
rect 2424 7954 2452 8298
rect 2412 7948 2464 7954
rect 2412 7890 2464 7896
rect 2792 7410 2820 9318
rect 2884 8906 2912 9454
rect 3056 9104 3108 9110
rect 3056 9046 3108 9052
rect 2872 8900 2924 8906
rect 2872 8842 2924 8848
rect 2884 8430 2912 8842
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 2964 7812 3016 7818
rect 2964 7754 3016 7760
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2976 7342 3004 7754
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 2504 7268 2556 7274
rect 2504 7210 2556 7216
rect 2516 6934 2544 7210
rect 2504 6928 2556 6934
rect 2504 6870 2556 6876
rect 2136 6860 2188 6866
rect 2136 6802 2188 6808
rect 2044 6792 2096 6798
rect 2044 6734 2096 6740
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 1584 6248 1636 6254
rect 1584 6190 1636 6196
rect 1858 6216 1914 6225
rect 1596 5166 1624 6190
rect 1858 6151 1914 6160
rect 1872 5914 1900 6151
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 2056 5710 2084 6734
rect 2148 6390 2176 6802
rect 2136 6384 2188 6390
rect 2136 6326 2188 6332
rect 2516 6254 2544 6870
rect 2780 6860 2832 6866
rect 2780 6802 2832 6808
rect 2504 6248 2556 6254
rect 2504 6190 2556 6196
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 1584 5160 1636 5166
rect 1584 5102 1636 5108
rect 480 4140 532 4146
rect 480 4082 532 4088
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 492 800 520 4082
rect 1492 3596 1544 3602
rect 1492 3538 1544 3544
rect 1400 2984 1452 2990
rect 1400 2926 1452 2932
rect 1412 800 1440 2926
rect 1504 2922 1532 3538
rect 1596 3058 1624 5102
rect 2136 5024 2188 5030
rect 2136 4966 2188 4972
rect 2148 4690 2176 4966
rect 2044 4684 2096 4690
rect 2044 4626 2096 4632
rect 2136 4684 2188 4690
rect 2136 4626 2188 4632
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 1964 4078 1992 4558
rect 2056 4214 2084 4626
rect 2044 4208 2096 4214
rect 2044 4150 2096 4156
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 1952 4072 2004 4078
rect 2136 4072 2188 4078
rect 1952 4014 2004 4020
rect 2056 4032 2136 4060
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 1584 3052 1636 3058
rect 1584 2994 1636 3000
rect 1688 2990 1716 3538
rect 1780 3466 1808 4014
rect 1860 3596 1912 3602
rect 1860 3538 1912 3544
rect 1768 3460 1820 3466
rect 1768 3402 1820 3408
rect 1676 2984 1728 2990
rect 1676 2926 1728 2932
rect 1492 2916 1544 2922
rect 1492 2858 1544 2864
rect 1872 2145 1900 3538
rect 1964 3126 1992 4014
rect 2056 3602 2084 4032
rect 2136 4014 2188 4020
rect 2228 3936 2280 3942
rect 2228 3878 2280 3884
rect 2240 3602 2268 3878
rect 2044 3596 2096 3602
rect 2044 3538 2096 3544
rect 2228 3596 2280 3602
rect 2228 3538 2280 3544
rect 1952 3120 2004 3126
rect 1952 3062 2004 3068
rect 1952 2916 2004 2922
rect 1952 2858 2004 2864
rect 1964 2514 1992 2858
rect 2504 2848 2556 2854
rect 2504 2790 2556 2796
rect 2516 2514 2544 2790
rect 1952 2508 2004 2514
rect 1952 2450 2004 2456
rect 2320 2508 2372 2514
rect 2320 2450 2372 2456
rect 2504 2508 2556 2514
rect 2504 2450 2556 2456
rect 1858 2136 1914 2145
rect 1858 2071 1914 2080
rect 1964 1426 1992 2450
rect 2332 2378 2360 2450
rect 2320 2372 2372 2378
rect 2320 2314 2372 2320
rect 2332 2106 2360 2314
rect 2320 2100 2372 2106
rect 2320 2042 2372 2048
rect 2686 1456 2742 1465
rect 1952 1420 2004 1426
rect 2686 1391 2688 1400
rect 1952 1362 2004 1368
rect 2740 1391 2742 1400
rect 2688 1362 2740 1368
rect 2792 800 2820 6802
rect 2872 6384 2924 6390
rect 2872 6326 2924 6332
rect 2884 5710 2912 6326
rect 3068 5846 3096 9046
rect 3056 5840 3108 5846
rect 3056 5782 3108 5788
rect 2872 5704 2924 5710
rect 2870 5672 2872 5681
rect 2924 5672 2926 5681
rect 2870 5607 2926 5616
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 2872 4480 2924 4486
rect 2872 4422 2924 4428
rect 2884 4282 2912 4422
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 2976 4078 3004 4558
rect 3252 4185 3280 9454
rect 3344 9110 3372 9658
rect 3514 9616 3570 9625
rect 3514 9551 3570 9560
rect 3528 9518 3556 9551
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 3608 9444 3660 9450
rect 3608 9386 3660 9392
rect 3332 9104 3384 9110
rect 3332 9046 3384 9052
rect 3332 8968 3384 8974
rect 3332 8910 3384 8916
rect 3344 8566 3372 8910
rect 3332 8560 3384 8566
rect 3332 8502 3384 8508
rect 3620 8430 3648 9386
rect 3608 8424 3660 8430
rect 3608 8366 3660 8372
rect 3896 8022 3924 13874
rect 4804 13864 4856 13870
rect 4908 13852 4936 14894
rect 4856 13824 4936 13852
rect 4804 13806 4856 13812
rect 4816 13462 4844 13806
rect 4804 13456 4856 13462
rect 4804 13398 4856 13404
rect 4712 13388 4764 13394
rect 4712 13330 4764 13336
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 4344 12912 4396 12918
rect 4344 12854 4396 12860
rect 4356 12442 4384 12854
rect 4724 12850 4752 13330
rect 5000 12866 5028 15574
rect 5816 15496 5868 15502
rect 5816 15438 5868 15444
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5460 14550 5488 15302
rect 5448 14544 5500 14550
rect 5448 14486 5500 14492
rect 5828 13870 5856 15438
rect 6012 15162 6040 16200
rect 6552 15564 6604 15570
rect 6552 15506 6604 15512
rect 6828 15564 6880 15570
rect 6828 15506 6880 15512
rect 6460 15496 6512 15502
rect 6460 15438 6512 15444
rect 6000 15156 6052 15162
rect 6000 15098 6052 15104
rect 6472 14482 6500 15438
rect 6564 14482 6592 15506
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6656 14958 6684 15302
rect 6644 14952 6696 14958
rect 6644 14894 6696 14900
rect 6736 14816 6788 14822
rect 6736 14758 6788 14764
rect 5908 14476 5960 14482
rect 5908 14418 5960 14424
rect 6460 14476 6512 14482
rect 6460 14418 6512 14424
rect 6552 14476 6604 14482
rect 6552 14418 6604 14424
rect 5920 14074 5948 14418
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 5816 13864 5868 13870
rect 5816 13806 5868 13812
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5356 13388 5408 13394
rect 5356 13330 5408 13336
rect 5172 13320 5224 13326
rect 5172 13262 5224 13268
rect 5080 13184 5132 13190
rect 5080 13126 5132 13132
rect 5092 12986 5120 13126
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 4712 12844 4764 12850
rect 5000 12838 5120 12866
rect 4712 12786 4764 12792
rect 4344 12436 4396 12442
rect 4724 12434 4752 12786
rect 4804 12708 4856 12714
rect 4804 12650 4856 12656
rect 4344 12378 4396 12384
rect 4632 12406 4752 12434
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 3976 11688 4028 11694
rect 3976 11630 4028 11636
rect 3988 11286 4016 11630
rect 4080 11626 4108 12242
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 4068 11620 4120 11626
rect 4068 11562 4120 11568
rect 3976 11280 4028 11286
rect 3976 11222 4028 11228
rect 4080 10538 4108 11562
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 4632 10742 4660 12406
rect 4816 12374 4844 12650
rect 4894 12472 4950 12481
rect 4894 12407 4950 12416
rect 4804 12368 4856 12374
rect 4804 12310 4856 12316
rect 4908 12170 4936 12407
rect 4896 12164 4948 12170
rect 4896 12106 4948 12112
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 4620 10736 4672 10742
rect 4620 10678 4672 10684
rect 4068 10532 4120 10538
rect 4068 10474 4120 10480
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3988 10305 4016 10406
rect 3974 10296 4030 10305
rect 3974 10231 4030 10240
rect 4632 10198 4660 10678
rect 4620 10192 4672 10198
rect 4620 10134 4672 10140
rect 3976 9988 4028 9994
rect 3976 9930 4028 9936
rect 4068 9988 4120 9994
rect 4068 9930 4120 9936
rect 3884 8016 3936 8022
rect 3884 7958 3936 7964
rect 3988 7954 4016 9930
rect 3332 7948 3384 7954
rect 3332 7890 3384 7896
rect 3976 7948 4028 7954
rect 3976 7890 4028 7896
rect 3344 7342 3372 7890
rect 3332 7336 3384 7342
rect 3332 7278 3384 7284
rect 3516 7336 3568 7342
rect 3516 7278 3568 7284
rect 3528 6662 3556 7278
rect 3792 7268 3844 7274
rect 3792 7210 3844 7216
rect 3804 6848 3832 7210
rect 4080 7002 4108 9930
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 4632 9518 4660 9862
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4724 9042 4752 11494
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 4160 8356 4212 8362
rect 4160 8298 4212 8304
rect 4172 8090 4200 8298
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 4344 7336 4396 7342
rect 4632 7290 4660 8910
rect 4344 7278 4396 7284
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 4356 6866 4384 7278
rect 4540 7274 4752 7290
rect 4528 7268 4752 7274
rect 4580 7262 4752 7268
rect 4528 7210 4580 7216
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 3884 6860 3936 6866
rect 3804 6820 3884 6848
rect 3884 6802 3936 6808
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3332 6180 3384 6186
rect 3332 6122 3384 6128
rect 3344 5778 3372 6122
rect 3528 5778 3556 6598
rect 3896 6322 3924 6802
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 3332 5772 3384 5778
rect 3332 5714 3384 5720
rect 3516 5772 3568 5778
rect 3516 5714 3568 5720
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 3608 5092 3660 5098
rect 3608 5034 3660 5040
rect 3620 4826 3648 5034
rect 3608 4820 3660 4826
rect 3608 4762 3660 4768
rect 3424 4684 3476 4690
rect 3424 4626 3476 4632
rect 3238 4176 3294 4185
rect 3238 4111 3294 4120
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 3332 4004 3384 4010
rect 3332 3946 3384 3952
rect 3056 3596 3108 3602
rect 3056 3538 3108 3544
rect 3068 2582 3096 3538
rect 3344 3534 3372 3946
rect 3436 3942 3464 4626
rect 3884 4616 3936 4622
rect 3884 4558 3936 4564
rect 3896 4078 3924 4558
rect 3884 4072 3936 4078
rect 3884 4014 3936 4020
rect 3896 3942 3924 4014
rect 3424 3936 3476 3942
rect 3424 3878 3476 3884
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3332 3528 3384 3534
rect 3332 3470 3384 3476
rect 4080 3058 4108 5102
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4172 4690 4200 4762
rect 4356 4690 4384 5170
rect 4632 5166 4660 7142
rect 4724 5778 4752 7262
rect 4816 5846 4844 11018
rect 4908 10130 4936 12106
rect 5092 11830 5120 12838
rect 5184 12306 5212 13262
rect 5368 12714 5396 13330
rect 5356 12708 5408 12714
rect 5408 12668 5488 12696
rect 5356 12650 5408 12656
rect 5264 12368 5316 12374
rect 5264 12310 5316 12316
rect 5172 12300 5224 12306
rect 5172 12242 5224 12248
rect 5184 12102 5212 12242
rect 5172 12096 5224 12102
rect 5172 12038 5224 12044
rect 5080 11824 5132 11830
rect 5080 11766 5132 11772
rect 5184 11218 5212 12038
rect 5276 11626 5304 12310
rect 5460 12306 5488 12668
rect 5552 12442 5580 13670
rect 5724 13388 5776 13394
rect 5724 13330 5776 13336
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5448 12300 5500 12306
rect 5448 12242 5500 12248
rect 5264 11620 5316 11626
rect 5264 11562 5316 11568
rect 5080 11212 5132 11218
rect 5080 11154 5132 11160
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 4988 10192 5040 10198
rect 4988 10134 5040 10140
rect 4896 10124 4948 10130
rect 4896 10066 4948 10072
rect 4896 9920 4948 9926
rect 4896 9862 4948 9868
rect 4908 9654 4936 9862
rect 4896 9648 4948 9654
rect 4896 9590 4948 9596
rect 5000 9178 5028 10134
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 4908 8294 4936 8978
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 5092 7274 5120 11154
rect 5184 10266 5212 11154
rect 5276 10674 5304 11562
rect 5356 11552 5408 11558
rect 5356 11494 5408 11500
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 5172 10260 5224 10266
rect 5172 10202 5224 10208
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 5184 9178 5212 10066
rect 5276 9518 5304 10610
rect 5368 10538 5396 11494
rect 5460 11218 5488 12242
rect 5632 12096 5684 12102
rect 5632 12038 5684 12044
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5448 10600 5500 10606
rect 5552 10588 5580 11698
rect 5644 11626 5672 12038
rect 5632 11620 5684 11626
rect 5632 11562 5684 11568
rect 5736 11558 5764 13330
rect 5828 12850 5856 13806
rect 6368 13456 6420 13462
rect 6368 13398 6420 13404
rect 5908 13388 5960 13394
rect 5908 13330 5960 13336
rect 5816 12844 5868 12850
rect 5816 12786 5868 12792
rect 5828 12481 5856 12786
rect 5814 12472 5870 12481
rect 5814 12407 5870 12416
rect 5920 11642 5948 13330
rect 6276 12708 6328 12714
rect 6276 12650 6328 12656
rect 6000 12640 6052 12646
rect 6000 12582 6052 12588
rect 6012 11898 6040 12582
rect 6288 12434 6316 12650
rect 6196 12406 6316 12434
rect 6092 12164 6144 12170
rect 6092 12106 6144 12112
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 6104 11762 6132 12106
rect 6092 11756 6144 11762
rect 6092 11698 6144 11704
rect 5920 11614 6040 11642
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5736 11200 5764 11494
rect 5920 11286 5948 11494
rect 5908 11280 5960 11286
rect 5908 11222 5960 11228
rect 5736 11172 5856 11200
rect 5724 11076 5776 11082
rect 5724 11018 5776 11024
rect 5500 10560 5580 10588
rect 5448 10542 5500 10548
rect 5356 10532 5408 10538
rect 5356 10474 5408 10480
rect 5368 10130 5396 10474
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5460 9926 5488 10202
rect 5448 9920 5500 9926
rect 5448 9862 5500 9868
rect 5264 9512 5316 9518
rect 5316 9472 5396 9500
rect 5264 9454 5316 9460
rect 5172 9172 5224 9178
rect 5172 9114 5224 9120
rect 5184 9042 5212 9114
rect 5264 9104 5316 9110
rect 5264 9046 5316 9052
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 5276 7410 5304 9046
rect 5368 8634 5396 9472
rect 5460 9382 5488 9862
rect 5552 9722 5580 10560
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 5540 9716 5592 9722
rect 5540 9658 5592 9664
rect 5644 9586 5672 9998
rect 5736 9722 5764 11018
rect 5828 11014 5856 11172
rect 5816 11008 5868 11014
rect 5816 10950 5868 10956
rect 5920 10690 5948 11222
rect 6012 11218 6040 11614
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 6012 10810 6040 11154
rect 6104 11150 6132 11698
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 5828 10662 5948 10690
rect 5828 10198 5856 10662
rect 5908 10600 5960 10606
rect 5908 10542 5960 10548
rect 5816 10192 5868 10198
rect 5816 10134 5868 10140
rect 5920 10130 5948 10542
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 5816 9920 5868 9926
rect 5816 9862 5868 9868
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5828 9450 5856 9862
rect 5632 9444 5684 9450
rect 5632 9386 5684 9392
rect 5816 9444 5868 9450
rect 5816 9386 5868 9392
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5460 8906 5488 9318
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5448 8900 5500 8906
rect 5448 8842 5500 8848
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5368 7954 5396 8570
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5080 7268 5132 7274
rect 5080 7210 5132 7216
rect 5460 6662 5488 7346
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5262 6352 5318 6361
rect 5460 6322 5488 6598
rect 5262 6287 5264 6296
rect 5316 6287 5318 6296
rect 5448 6316 5500 6322
rect 5264 6258 5316 6264
rect 5448 6258 5500 6264
rect 5552 6254 5580 9114
rect 5644 8922 5672 9386
rect 5644 8906 5764 8922
rect 5644 8900 5776 8906
rect 5644 8894 5724 8900
rect 5724 8842 5776 8848
rect 5816 8424 5868 8430
rect 5816 8366 5868 8372
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 5644 8090 5672 8298
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 5828 7954 5856 8366
rect 5920 8294 5948 10066
rect 6104 9926 6132 11086
rect 6092 9920 6144 9926
rect 6092 9862 6144 9868
rect 6092 9104 6144 9110
rect 6092 9046 6144 9052
rect 6104 8634 6132 9046
rect 6196 8650 6224 12406
rect 6380 12102 6408 13398
rect 6472 13394 6500 14418
rect 6564 13462 6592 14418
rect 6748 14414 6776 14758
rect 6736 14408 6788 14414
rect 6736 14350 6788 14356
rect 6840 14346 6868 15506
rect 6932 15026 6960 16200
rect 8312 15994 8340 16200
rect 8312 15966 8616 15994
rect 8220 15804 8516 15824
rect 8276 15802 8300 15804
rect 8356 15802 8380 15804
rect 8436 15802 8460 15804
rect 8298 15750 8300 15802
rect 8362 15750 8374 15802
rect 8436 15750 8438 15802
rect 8276 15748 8300 15750
rect 8356 15748 8380 15750
rect 8436 15748 8460 15750
rect 8220 15728 8516 15748
rect 8588 15586 8616 15966
rect 8496 15558 8616 15586
rect 8760 15564 8812 15570
rect 8024 15496 8076 15502
rect 8024 15438 8076 15444
rect 7012 15428 7064 15434
rect 7012 15370 7064 15376
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 6828 14340 6880 14346
rect 6828 14282 6880 14288
rect 6840 14006 6868 14282
rect 6828 14000 6880 14006
rect 6828 13942 6880 13948
rect 7024 13938 7052 15370
rect 7288 15360 7340 15366
rect 7288 15302 7340 15308
rect 7300 14550 7328 15302
rect 7932 15020 7984 15026
rect 7932 14962 7984 14968
rect 7288 14544 7340 14550
rect 7288 14486 7340 14492
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 7012 13932 7064 13938
rect 7012 13874 7064 13880
rect 7576 13870 7604 14418
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 6552 13456 6604 13462
rect 6552 13398 6604 13404
rect 6460 13388 6512 13394
rect 6460 13330 6512 13336
rect 7380 13252 7432 13258
rect 7380 13194 7432 13200
rect 6828 13184 6880 13190
rect 6828 13126 6880 13132
rect 6552 12912 6604 12918
rect 6552 12854 6604 12860
rect 6368 12096 6420 12102
rect 6368 12038 6420 12044
rect 6380 11626 6408 12038
rect 6564 11898 6592 12854
rect 6840 12238 6868 13126
rect 6920 12708 6972 12714
rect 6920 12650 6972 12656
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 6932 12186 6960 12650
rect 7392 12646 7420 13194
rect 7576 12986 7604 13806
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7472 12776 7524 12782
rect 7472 12718 7524 12724
rect 7012 12640 7064 12646
rect 7012 12582 7064 12588
rect 7380 12640 7432 12646
rect 7380 12582 7432 12588
rect 7024 12442 7052 12582
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6460 11688 6512 11694
rect 6460 11630 6512 11636
rect 6368 11620 6420 11626
rect 6368 11562 6420 11568
rect 6380 10062 6408 11562
rect 6472 11218 6500 11630
rect 6460 11212 6512 11218
rect 6460 11154 6512 11160
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 6092 8628 6144 8634
rect 6196 8622 6316 8650
rect 6092 8570 6144 8576
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 6196 8090 6224 8434
rect 6184 8084 6236 8090
rect 6184 8026 6236 8032
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5632 7268 5684 7274
rect 5632 7210 5684 7216
rect 5644 6866 5672 7210
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5828 6730 5856 7482
rect 5816 6724 5868 6730
rect 5816 6666 5868 6672
rect 5920 6390 5948 7686
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 5816 6384 5868 6390
rect 5816 6326 5868 6332
rect 5908 6384 5960 6390
rect 5908 6326 5960 6332
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 4804 5840 4856 5846
rect 4804 5782 4856 5788
rect 4712 5772 4764 5778
rect 4712 5714 4764 5720
rect 5632 5772 5684 5778
rect 5632 5714 5684 5720
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 5356 4752 5408 4758
rect 5356 4694 5408 4700
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 4620 4548 4672 4554
rect 4620 4490 4672 4496
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 4436 4208 4488 4214
rect 4436 4150 4488 4156
rect 4448 3534 4476 4150
rect 4632 4026 4660 4490
rect 4540 3998 4660 4026
rect 4540 3602 4568 3998
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 4632 3670 4660 3878
rect 4620 3664 4672 3670
rect 4620 3606 4672 3612
rect 4528 3596 4580 3602
rect 4528 3538 4580 3544
rect 4436 3528 4488 3534
rect 4436 3470 4488 3476
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 4632 3194 4660 3606
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4724 3074 4752 3878
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 4632 3046 4752 3074
rect 3792 2916 3844 2922
rect 3792 2858 3844 2864
rect 3424 2848 3476 2854
rect 3424 2790 3476 2796
rect 3056 2576 3108 2582
rect 3056 2518 3108 2524
rect 3332 2508 3384 2514
rect 3436 2496 3464 2790
rect 3384 2468 3464 2496
rect 3332 2450 3384 2456
rect 3804 2378 3832 2858
rect 3332 2372 3384 2378
rect 3332 2314 3384 2320
rect 3792 2372 3844 2378
rect 3792 2314 3844 2320
rect 2872 1828 2924 1834
rect 2872 1770 2924 1776
rect 2884 1562 2912 1770
rect 2872 1556 2924 1562
rect 2872 1498 2924 1504
rect 3344 1426 3372 2314
rect 4080 1970 4108 2994
rect 4632 2650 4660 3046
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4160 2508 4212 2514
rect 4160 2450 4212 2456
rect 4172 2378 4200 2450
rect 4724 2394 4752 2926
rect 4804 2848 4856 2854
rect 4804 2790 4856 2796
rect 4816 2582 4844 2790
rect 4804 2576 4856 2582
rect 4804 2518 4856 2524
rect 4632 2378 4752 2394
rect 4160 2372 4212 2378
rect 4160 2314 4212 2320
rect 4620 2372 4752 2378
rect 4672 2366 4752 2372
rect 4620 2314 4672 2320
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 4632 2106 4660 2314
rect 4620 2100 4672 2106
rect 4620 2042 4672 2048
rect 4252 2032 4304 2038
rect 4252 1974 4304 1980
rect 4068 1964 4120 1970
rect 4068 1906 4120 1912
rect 4160 1964 4212 1970
rect 4160 1906 4212 1912
rect 3976 1760 4028 1766
rect 3976 1702 4028 1708
rect 3988 1426 4016 1702
rect 3332 1420 3384 1426
rect 3332 1362 3384 1368
rect 3976 1420 4028 1426
rect 3976 1362 4028 1368
rect 4080 1222 4108 1906
rect 4172 1290 4200 1906
rect 4264 1426 4292 1974
rect 4632 1902 4660 2042
rect 4908 1986 4936 4558
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 4816 1970 4936 1986
rect 4804 1964 4936 1970
rect 4856 1958 4936 1964
rect 4804 1906 4856 1912
rect 4620 1896 4672 1902
rect 4620 1838 4672 1844
rect 4620 1760 4672 1766
rect 4620 1702 4672 1708
rect 4252 1420 4304 1426
rect 4252 1362 4304 1368
rect 4632 1358 4660 1702
rect 4620 1352 4672 1358
rect 4620 1294 4672 1300
rect 4160 1284 4212 1290
rect 4160 1226 4212 1232
rect 4068 1216 4120 1222
rect 4068 1158 4120 1164
rect 4220 1116 4516 1136
rect 4276 1114 4300 1116
rect 4356 1114 4380 1116
rect 4436 1114 4460 1116
rect 4298 1062 4300 1114
rect 4362 1062 4374 1114
rect 4436 1062 4438 1114
rect 4276 1060 4300 1062
rect 4356 1060 4380 1062
rect 4436 1060 4460 1062
rect 4220 1040 4516 1060
rect 5000 898 5028 3878
rect 5368 3738 5396 4694
rect 5552 4554 5580 5510
rect 5644 5370 5672 5714
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5828 5098 5856 6326
rect 6196 5846 6224 6802
rect 6184 5840 6236 5846
rect 6184 5782 6236 5788
rect 6000 5364 6052 5370
rect 6000 5306 6052 5312
rect 6012 5166 6040 5306
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 5724 5092 5776 5098
rect 5724 5034 5776 5040
rect 5816 5092 5868 5098
rect 5816 5034 5868 5040
rect 5736 4826 5764 5034
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 5540 4548 5592 4554
rect 5540 4490 5592 4496
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 5644 3738 5672 3946
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5368 2650 5396 3674
rect 5460 3398 5488 3674
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 5368 2514 5396 2586
rect 5172 2508 5224 2514
rect 5172 2450 5224 2456
rect 5356 2508 5408 2514
rect 5356 2450 5408 2456
rect 5184 1834 5212 2450
rect 5368 2310 5396 2450
rect 5356 2304 5408 2310
rect 5356 2246 5408 2252
rect 5368 1902 5396 2246
rect 5460 2038 5488 3334
rect 5552 3126 5580 3538
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 5644 3126 5672 3470
rect 5540 3120 5592 3126
rect 5540 3062 5592 3068
rect 5632 3120 5684 3126
rect 5632 3062 5684 3068
rect 5644 2650 5672 3062
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 5448 2032 5500 2038
rect 5448 1974 5500 1980
rect 5356 1896 5408 1902
rect 5356 1838 5408 1844
rect 5172 1828 5224 1834
rect 5172 1770 5224 1776
rect 4172 870 5028 898
rect 4172 800 4200 870
rect 5552 800 5580 2246
rect 5644 1902 5672 2450
rect 5736 2378 5764 4558
rect 6012 4078 6040 5102
rect 6000 4072 6052 4078
rect 6000 4014 6052 4020
rect 5908 3596 5960 3602
rect 5908 3538 5960 3544
rect 5816 3460 5868 3466
rect 5816 3402 5868 3408
rect 5828 2854 5856 3402
rect 5920 2990 5948 3538
rect 5908 2984 5960 2990
rect 5908 2926 5960 2932
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 5828 2378 5856 2790
rect 6012 2774 6040 4014
rect 6288 3942 6316 8622
rect 6368 7812 6420 7818
rect 6368 7754 6420 7760
rect 6380 5846 6408 7754
rect 6472 6866 6500 11154
rect 6564 10169 6592 11834
rect 6736 11824 6788 11830
rect 6736 11766 6788 11772
rect 6748 11218 6776 11766
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6748 10538 6776 11154
rect 6840 11082 6868 12174
rect 6932 12158 7144 12186
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 6932 11150 6960 12038
rect 7024 11218 7052 12038
rect 7012 11212 7064 11218
rect 7012 11154 7064 11160
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 6828 11076 6880 11082
rect 6828 11018 6880 11024
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 6736 10532 6788 10538
rect 6736 10474 6788 10480
rect 6748 10266 6776 10474
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 6550 10160 6606 10169
rect 6550 10095 6552 10104
rect 6604 10095 6606 10104
rect 6552 10066 6604 10072
rect 6564 10035 6592 10066
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6564 7342 6592 8230
rect 6656 8090 6684 9998
rect 6840 9674 6868 10746
rect 6932 10130 6960 11086
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 7024 9722 7052 10610
rect 7116 10470 7144 12158
rect 7208 11218 7236 12378
rect 7484 12356 7512 12718
rect 7564 12368 7616 12374
rect 7484 12328 7564 12356
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7288 12164 7340 12170
rect 7288 12106 7340 12112
rect 7300 11762 7328 12106
rect 7288 11756 7340 11762
rect 7288 11698 7340 11704
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 7300 10606 7328 11698
rect 7392 11694 7420 12242
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7484 10674 7512 12328
rect 7564 12310 7616 12316
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 6748 9654 6868 9674
rect 7012 9716 7064 9722
rect 7012 9658 7064 9664
rect 6748 9648 6880 9654
rect 6748 9646 6828 9648
rect 6748 8838 6776 9646
rect 6828 9590 6880 9596
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 6840 8430 6868 9114
rect 7024 8498 7052 9318
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7116 8634 7144 8774
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 7300 8362 7328 10542
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 7392 9450 7420 9862
rect 7380 9444 7432 9450
rect 7380 9386 7432 9392
rect 7472 9444 7524 9450
rect 7472 9386 7524 9392
rect 7288 8356 7340 8362
rect 7288 8298 7340 8304
rect 6644 8084 6696 8090
rect 6644 8026 6696 8032
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 7196 7948 7248 7954
rect 7196 7890 7248 7896
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6840 7478 6868 7822
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 6736 7268 6788 7274
rect 6736 7210 6788 7216
rect 6460 6860 6512 6866
rect 6460 6802 6512 6808
rect 6748 5914 6776 7210
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6368 5840 6420 5846
rect 6368 5782 6420 5788
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6380 4690 6408 4966
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6380 4010 6408 4626
rect 6368 4004 6420 4010
rect 6368 3946 6420 3952
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 6276 2984 6328 2990
rect 6276 2926 6328 2932
rect 6012 2746 6224 2774
rect 6196 2514 6224 2746
rect 6288 2582 6316 2926
rect 6380 2650 6408 3946
rect 6564 3602 6592 4966
rect 6736 4752 6788 4758
rect 6736 4694 6788 4700
rect 6748 4078 6776 4694
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 6840 4010 6868 4626
rect 6828 4004 6880 4010
rect 6828 3946 6880 3952
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 6564 3194 6592 3538
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 6748 2990 6776 3878
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 6276 2576 6328 2582
rect 6276 2518 6328 2524
rect 6184 2508 6236 2514
rect 6184 2450 6236 2456
rect 5724 2372 5776 2378
rect 5724 2314 5776 2320
rect 5816 2372 5868 2378
rect 5816 2314 5868 2320
rect 5632 1896 5684 1902
rect 5632 1838 5684 1844
rect 5736 1850 5764 2314
rect 5828 1970 5856 2314
rect 5816 1964 5868 1970
rect 5816 1906 5868 1912
rect 6000 1896 6052 1902
rect 5736 1844 6000 1850
rect 5736 1838 6052 1844
rect 5736 1822 6040 1838
rect 6196 1766 6224 2450
rect 6288 2106 6316 2518
rect 6552 2508 6604 2514
rect 6552 2450 6604 2456
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 6276 2100 6328 2106
rect 6276 2042 6328 2048
rect 6564 1902 6592 2450
rect 6644 2372 6696 2378
rect 6644 2314 6696 2320
rect 6552 1896 6604 1902
rect 6552 1838 6604 1844
rect 6184 1760 6236 1766
rect 6184 1702 6236 1708
rect 6196 1222 6224 1702
rect 6656 1562 6684 2314
rect 6748 1562 6776 2450
rect 6828 1760 6880 1766
rect 6828 1702 6880 1708
rect 6644 1556 6696 1562
rect 6644 1498 6696 1504
rect 6736 1556 6788 1562
rect 6736 1498 6788 1504
rect 6840 1358 6868 1702
rect 6828 1352 6880 1358
rect 6828 1294 6880 1300
rect 6184 1216 6236 1222
rect 6184 1158 6236 1164
rect 6932 800 6960 7890
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 7024 6254 7052 6938
rect 7208 6662 7236 7890
rect 7300 7750 7328 8298
rect 7392 7954 7420 9386
rect 7484 9110 7512 9386
rect 7472 9104 7524 9110
rect 7472 9046 7524 9052
rect 7564 9036 7616 9042
rect 7564 8978 7616 8984
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7300 6254 7328 7686
rect 7380 7268 7432 7274
rect 7380 7210 7432 7216
rect 7392 6662 7420 7210
rect 7484 6934 7512 8910
rect 7576 8430 7604 8978
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7472 6928 7524 6934
rect 7472 6870 7524 6876
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7012 6248 7064 6254
rect 7012 6190 7064 6196
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7288 6248 7340 6254
rect 7288 6190 7340 6196
rect 7208 5846 7236 6190
rect 7196 5840 7248 5846
rect 7196 5782 7248 5788
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 7392 4690 7420 5510
rect 7484 5370 7512 6870
rect 7576 6390 7604 8366
rect 7668 7546 7696 13330
rect 7944 13326 7972 14962
rect 8036 14958 8064 15438
rect 8496 15026 8524 15558
rect 8760 15506 8812 15512
rect 8576 15360 8628 15366
rect 8576 15302 8628 15308
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8024 14952 8076 14958
rect 8024 14894 8076 14900
rect 8588 14890 8616 15302
rect 8772 14890 8800 15506
rect 9692 14906 9720 16200
rect 10232 15564 10284 15570
rect 10232 15506 10284 15512
rect 10140 15360 10192 15366
rect 10140 15302 10192 15308
rect 9862 15056 9918 15065
rect 9862 14991 9864 15000
rect 9916 14991 9918 15000
rect 9864 14962 9916 14968
rect 8576 14884 8628 14890
rect 8576 14826 8628 14832
rect 8760 14884 8812 14890
rect 9692 14878 9904 14906
rect 8760 14826 8812 14832
rect 8024 14816 8076 14822
rect 8024 14758 8076 14764
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 7760 12306 7788 12718
rect 7944 12714 7972 13262
rect 8036 12986 8064 14758
rect 8220 14716 8516 14736
rect 8276 14714 8300 14716
rect 8356 14714 8380 14716
rect 8436 14714 8460 14716
rect 8298 14662 8300 14714
rect 8362 14662 8374 14714
rect 8436 14662 8438 14714
rect 8276 14660 8300 14662
rect 8356 14660 8380 14662
rect 8436 14660 8460 14662
rect 8220 14640 8516 14660
rect 8588 14618 8616 14826
rect 8576 14612 8628 14618
rect 8576 14554 8628 14560
rect 8668 14340 8720 14346
rect 8668 14282 8720 14288
rect 8680 14074 8708 14282
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8576 14000 8628 14006
rect 8576 13942 8628 13948
rect 8220 13628 8516 13648
rect 8276 13626 8300 13628
rect 8356 13626 8380 13628
rect 8436 13626 8460 13628
rect 8298 13574 8300 13626
rect 8362 13574 8374 13626
rect 8436 13574 8438 13626
rect 8276 13572 8300 13574
rect 8356 13572 8380 13574
rect 8436 13572 8460 13574
rect 8220 13552 8516 13572
rect 8588 13462 8616 13942
rect 8772 13870 8800 14826
rect 9220 14816 9272 14822
rect 9220 14758 9272 14764
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 9232 14482 9260 14758
rect 8852 14476 8904 14482
rect 8852 14418 8904 14424
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8772 13462 8800 13806
rect 8864 13530 8892 14418
rect 9232 13938 9260 14418
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 9312 13524 9364 13530
rect 9312 13466 9364 13472
rect 8576 13456 8628 13462
rect 8576 13398 8628 13404
rect 8760 13456 8812 13462
rect 8760 13398 8812 13404
rect 8116 13388 8168 13394
rect 8116 13330 8168 13336
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 7932 12708 7984 12714
rect 7932 12650 7984 12656
rect 8024 12708 8076 12714
rect 8024 12650 8076 12656
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 7840 11280 7892 11286
rect 7840 11222 7892 11228
rect 7852 10810 7880 11222
rect 7944 11218 7972 12650
rect 8036 12306 8064 12650
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 8128 12238 8156 13330
rect 8852 13320 8904 13326
rect 8852 13262 8904 13268
rect 8864 12850 8892 13262
rect 8944 12980 8996 12986
rect 8944 12922 8996 12928
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8668 12708 8720 12714
rect 8668 12650 8720 12656
rect 8852 12708 8904 12714
rect 8852 12650 8904 12656
rect 8576 12640 8628 12646
rect 8576 12582 8628 12588
rect 8220 12540 8516 12560
rect 8276 12538 8300 12540
rect 8356 12538 8380 12540
rect 8436 12538 8460 12540
rect 8298 12486 8300 12538
rect 8362 12486 8374 12538
rect 8436 12486 8438 12538
rect 8276 12484 8300 12486
rect 8356 12484 8380 12486
rect 8436 12484 8460 12486
rect 8220 12464 8516 12484
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 8392 12232 8444 12238
rect 8496 12209 8524 12242
rect 8392 12174 8444 12180
rect 8482 12200 8538 12209
rect 8404 11762 8432 12174
rect 8482 12135 8538 12144
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8496 11898 8524 12038
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8024 11688 8076 11694
rect 8496 11665 8524 11834
rect 8588 11830 8616 12582
rect 8576 11824 8628 11830
rect 8576 11766 8628 11772
rect 8024 11630 8076 11636
rect 8482 11656 8538 11665
rect 8036 11354 8064 11630
rect 8116 11620 8168 11626
rect 8482 11591 8538 11600
rect 8116 11562 8168 11568
rect 8024 11348 8076 11354
rect 8024 11290 8076 11296
rect 7932 11212 7984 11218
rect 7932 11154 7984 11160
rect 7840 10804 7892 10810
rect 7840 10746 7892 10752
rect 7840 10532 7892 10538
rect 7840 10474 7892 10480
rect 7932 10532 7984 10538
rect 7932 10474 7984 10480
rect 7748 10464 7800 10470
rect 7748 10406 7800 10412
rect 7760 10130 7788 10406
rect 7748 10124 7800 10130
rect 7748 10066 7800 10072
rect 7852 9994 7880 10474
rect 7840 9988 7892 9994
rect 7840 9930 7892 9936
rect 7944 9518 7972 10474
rect 8022 10160 8078 10169
rect 8128 10130 8156 11562
rect 8220 11452 8516 11472
rect 8276 11450 8300 11452
rect 8356 11450 8380 11452
rect 8436 11450 8460 11452
rect 8298 11398 8300 11450
rect 8362 11398 8374 11450
rect 8436 11398 8438 11450
rect 8276 11396 8300 11398
rect 8356 11396 8380 11398
rect 8436 11396 8460 11398
rect 8220 11376 8516 11396
rect 8220 10364 8516 10384
rect 8276 10362 8300 10364
rect 8356 10362 8380 10364
rect 8436 10362 8460 10364
rect 8298 10310 8300 10362
rect 8362 10310 8374 10362
rect 8436 10310 8438 10362
rect 8276 10308 8300 10310
rect 8356 10308 8380 10310
rect 8436 10308 8460 10310
rect 8220 10288 8516 10308
rect 8588 10130 8616 11766
rect 8680 11694 8708 12650
rect 8760 12300 8812 12306
rect 8760 12242 8812 12248
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8680 11218 8708 11494
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 8772 10266 8800 12242
rect 8864 11762 8892 12650
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8852 11144 8904 11150
rect 8852 11086 8904 11092
rect 8864 10606 8892 11086
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8022 10095 8024 10104
rect 8076 10095 8078 10104
rect 8116 10124 8168 10130
rect 8024 10066 8076 10072
rect 8116 10066 8168 10072
rect 8576 10124 8628 10130
rect 8576 10066 8628 10072
rect 8668 10124 8720 10130
rect 8668 10066 8720 10072
rect 8576 9988 8628 9994
rect 8576 9930 8628 9936
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 8022 9480 8078 9489
rect 8022 9415 8078 9424
rect 8116 9444 8168 9450
rect 7932 9376 7984 9382
rect 8036 9364 8064 9415
rect 8116 9386 8168 9392
rect 7984 9336 8064 9364
rect 7932 9318 7984 9324
rect 7840 8900 7892 8906
rect 7840 8842 7892 8848
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 7760 8022 7788 8366
rect 7748 8016 7800 8022
rect 7748 7958 7800 7964
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 7654 7440 7710 7449
rect 7654 7375 7710 7384
rect 7668 7274 7696 7375
rect 7656 7268 7708 7274
rect 7656 7210 7708 7216
rect 7668 6390 7696 7210
rect 7564 6384 7616 6390
rect 7564 6326 7616 6332
rect 7656 6384 7708 6390
rect 7656 6326 7708 6332
rect 7760 6118 7788 7958
rect 7852 7886 7880 8842
rect 7932 8560 7984 8566
rect 7932 8502 7984 8508
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7852 7002 7880 7822
rect 7840 6996 7892 7002
rect 7840 6938 7892 6944
rect 7944 6390 7972 8502
rect 8036 7857 8064 9336
rect 8128 8838 8156 9386
rect 8220 9276 8516 9296
rect 8276 9274 8300 9276
rect 8356 9274 8380 9276
rect 8436 9274 8460 9276
rect 8298 9222 8300 9274
rect 8362 9222 8374 9274
rect 8436 9222 8438 9274
rect 8276 9220 8300 9222
rect 8356 9220 8380 9222
rect 8436 9220 8460 9222
rect 8220 9200 8516 9220
rect 8588 9042 8616 9930
rect 8680 9450 8708 10066
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 8668 9444 8720 9450
rect 8668 9386 8720 9392
rect 8576 9036 8628 9042
rect 8576 8978 8628 8984
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 8220 8566 8248 8910
rect 8680 8634 8708 9386
rect 8772 9110 8800 9998
rect 8956 9738 8984 12922
rect 9220 12640 9272 12646
rect 9220 12582 9272 12588
rect 9128 12436 9180 12442
rect 9232 12424 9260 12582
rect 9324 12442 9352 13466
rect 9496 13388 9548 13394
rect 9496 13330 9548 13336
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9180 12396 9260 12424
rect 9128 12378 9180 12384
rect 9232 12084 9260 12396
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 9508 12374 9536 13330
rect 9692 12986 9720 13330
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9496 12368 9548 12374
rect 9496 12310 9548 12316
rect 9312 12096 9364 12102
rect 9232 12056 9312 12084
rect 9312 12038 9364 12044
rect 9220 11824 9272 11830
rect 9220 11766 9272 11772
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 9036 11280 9088 11286
rect 9036 11222 9088 11228
rect 8864 9710 8984 9738
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8760 8900 8812 8906
rect 8760 8842 8812 8848
rect 8772 8634 8800 8842
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8208 8560 8260 8566
rect 8208 8502 8260 8508
rect 8772 8430 8800 8570
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 8116 8356 8168 8362
rect 8116 8298 8168 8304
rect 8128 7954 8156 8298
rect 8220 8188 8516 8208
rect 8276 8186 8300 8188
rect 8356 8186 8380 8188
rect 8436 8186 8460 8188
rect 8298 8134 8300 8186
rect 8362 8134 8374 8186
rect 8436 8134 8438 8186
rect 8276 8132 8300 8134
rect 8356 8132 8380 8134
rect 8436 8132 8460 8134
rect 8220 8112 8516 8132
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 8022 7848 8078 7857
rect 8022 7783 8078 7792
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 7932 6384 7984 6390
rect 7932 6326 7984 6332
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 7852 5710 7880 6190
rect 7944 5846 7972 6326
rect 8036 6254 8064 7686
rect 8128 7478 8156 7890
rect 8116 7472 8168 7478
rect 8116 7414 8168 7420
rect 8208 7472 8260 7478
rect 8208 7414 8260 7420
rect 8220 7188 8248 7414
rect 8128 7160 8248 7188
rect 8668 7200 8720 7206
rect 8128 6458 8156 7160
rect 8668 7142 8720 7148
rect 8760 7200 8812 7206
rect 8760 7142 8812 7148
rect 8220 7100 8516 7120
rect 8276 7098 8300 7100
rect 8356 7098 8380 7100
rect 8436 7098 8460 7100
rect 8298 7046 8300 7098
rect 8362 7046 8374 7098
rect 8436 7046 8438 7098
rect 8276 7044 8300 7046
rect 8356 7044 8380 7046
rect 8436 7044 8460 7046
rect 8220 7024 8516 7044
rect 8680 6882 8708 7142
rect 8772 7002 8800 7142
rect 8760 6996 8812 7002
rect 8760 6938 8812 6944
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8496 6854 8708 6882
rect 8760 6860 8812 6866
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8220 6390 8248 6802
rect 8496 6730 8524 6854
rect 8760 6802 8812 6808
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 8484 6724 8536 6730
rect 8484 6666 8536 6672
rect 8208 6384 8260 6390
rect 8208 6326 8260 6332
rect 8680 6254 8708 6734
rect 8024 6248 8076 6254
rect 8024 6190 8076 6196
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8220 6012 8516 6032
rect 8276 6010 8300 6012
rect 8356 6010 8380 6012
rect 8436 6010 8460 6012
rect 8298 5958 8300 6010
rect 8362 5958 8374 6010
rect 8436 5958 8438 6010
rect 8276 5956 8300 5958
rect 8356 5956 8380 5958
rect 8436 5956 8460 5958
rect 8220 5936 8516 5956
rect 7932 5840 7984 5846
rect 7932 5782 7984 5788
rect 8772 5778 8800 6802
rect 8760 5772 8812 5778
rect 8760 5714 8812 5720
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8024 5568 8076 5574
rect 8484 5568 8536 5574
rect 8024 5510 8076 5516
rect 8482 5536 8484 5545
rect 8536 5536 8538 5545
rect 7472 5364 7524 5370
rect 7472 5306 7524 5312
rect 8036 5234 8064 5510
rect 8482 5471 8538 5480
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 8220 4924 8516 4944
rect 8276 4922 8300 4924
rect 8356 4922 8380 4924
rect 8436 4922 8460 4924
rect 8298 4870 8300 4922
rect 8362 4870 8374 4922
rect 8436 4870 8438 4922
rect 8276 4868 8300 4870
rect 8356 4868 8380 4870
rect 8436 4868 8460 4870
rect 8220 4848 8516 4868
rect 8680 4690 8708 5646
rect 8772 5370 8800 5714
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7656 4684 7708 4690
rect 7656 4626 7708 4632
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 7024 4010 7052 4558
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7392 4078 7420 4422
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 7380 4072 7432 4078
rect 7380 4014 7432 4020
rect 7012 4004 7064 4010
rect 7012 3946 7064 3952
rect 7024 3670 7052 3946
rect 7012 3664 7064 3670
rect 7012 3606 7064 3612
rect 7116 3602 7144 4014
rect 7668 3652 7696 4626
rect 8772 4622 8800 5306
rect 8864 4826 8892 9710
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 8956 8906 8984 9590
rect 8944 8900 8996 8906
rect 8944 8842 8996 8848
rect 8956 8430 8984 8842
rect 8944 8424 8996 8430
rect 8944 8366 8996 8372
rect 9048 7426 9076 11222
rect 9140 11082 9168 11698
rect 9232 11665 9260 11766
rect 9324 11694 9352 12038
rect 9680 11756 9732 11762
rect 9508 11716 9680 11744
rect 9312 11688 9364 11694
rect 9218 11656 9274 11665
rect 9508 11642 9536 11716
rect 9680 11698 9732 11704
rect 9312 11630 9364 11636
rect 9416 11626 9536 11642
rect 9218 11591 9274 11600
rect 9404 11620 9536 11626
rect 9456 11614 9536 11620
rect 9586 11656 9642 11665
rect 9586 11591 9642 11600
rect 9404 11562 9456 11568
rect 9402 11384 9458 11393
rect 9402 11319 9458 11328
rect 9128 11076 9180 11082
rect 9128 11018 9180 11024
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 9232 10538 9260 10950
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 9220 10532 9272 10538
rect 9220 10474 9272 10480
rect 9324 10130 9352 10542
rect 9312 10124 9364 10130
rect 9312 10066 9364 10072
rect 9220 9716 9272 9722
rect 9220 9658 9272 9664
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 9140 9194 9168 9590
rect 9232 9518 9260 9658
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 9324 9450 9352 10066
rect 9312 9444 9364 9450
rect 9312 9386 9364 9392
rect 9140 9166 9352 9194
rect 9220 9036 9272 9042
rect 9220 8978 9272 8984
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 9140 7954 9168 8774
rect 9232 8566 9260 8978
rect 9220 8560 9272 8566
rect 9220 8502 9272 8508
rect 9324 8498 9352 9166
rect 9416 9110 9444 11319
rect 9600 10810 9628 11591
rect 9784 11354 9812 14758
rect 9876 12850 9904 14878
rect 9956 14272 10008 14278
rect 9956 14214 10008 14220
rect 9968 14006 9996 14214
rect 9956 14000 10008 14006
rect 9956 13942 10008 13948
rect 10152 13938 10180 15302
rect 10244 14006 10272 15506
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10232 14000 10284 14006
rect 10232 13942 10284 13948
rect 10140 13932 10192 13938
rect 10140 13874 10192 13880
rect 10244 13462 10272 13942
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 10232 13456 10284 13462
rect 10232 13398 10284 13404
rect 10336 13394 10364 13806
rect 10324 13388 10376 13394
rect 10324 13330 10376 13336
rect 10428 13326 10456 15098
rect 10968 14476 11020 14482
rect 10968 14418 11020 14424
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 10888 13938 10916 14214
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 10980 13870 11008 14418
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 10980 13462 11008 13806
rect 10968 13456 11020 13462
rect 10968 13398 11020 13404
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 10232 12844 10286 12889
rect 10428 12850 10456 13262
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 10876 12912 10928 12918
rect 10876 12854 10928 12860
rect 10416 12844 10468 12850
rect 10232 12786 10284 12792
rect 10416 12786 10468 12792
rect 10324 12436 10376 12442
rect 10324 12378 10376 12384
rect 10232 12368 10284 12374
rect 10232 12310 10284 12316
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 9862 12200 9918 12209
rect 9862 12135 9918 12144
rect 9876 11558 9904 12135
rect 10152 11898 10180 12242
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10244 11626 10272 12310
rect 10232 11620 10284 11626
rect 10232 11562 10284 11568
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9876 11200 9904 11494
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 9956 11212 10008 11218
rect 9876 11172 9956 11200
rect 9956 11154 10008 11160
rect 9864 11008 9916 11014
rect 9864 10950 9916 10956
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 9876 10606 9904 10950
rect 9968 10674 9996 11154
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 9864 10600 9916 10606
rect 9784 10548 9864 10554
rect 9784 10542 9916 10548
rect 9784 10526 9904 10542
rect 9784 10130 9812 10526
rect 9956 10464 10008 10470
rect 10060 10452 10088 11222
rect 10232 10668 10284 10674
rect 10232 10610 10284 10616
rect 10008 10424 10088 10452
rect 9956 10406 10008 10412
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9508 9518 9536 10066
rect 9784 9674 9812 10066
rect 9692 9646 9812 9674
rect 9496 9512 9548 9518
rect 9692 9500 9720 9646
rect 9496 9454 9548 9460
rect 9586 9480 9642 9489
rect 9508 9178 9536 9454
rect 9692 9472 9812 9500
rect 9642 9424 9720 9432
rect 9586 9415 9720 9424
rect 9600 9404 9720 9415
rect 9692 9353 9720 9404
rect 9678 9344 9734 9353
rect 9678 9279 9734 9288
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9404 9104 9456 9110
rect 9404 9046 9456 9052
rect 9600 9024 9628 9114
rect 9508 8996 9628 9024
rect 9508 8838 9536 8996
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9692 8537 9720 8774
rect 9678 8528 9734 8537
rect 9312 8492 9364 8498
rect 9678 8463 9734 8472
rect 9312 8434 9364 8440
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9404 8356 9456 8362
rect 9404 8298 9456 8304
rect 9128 7948 9180 7954
rect 9128 7890 9180 7896
rect 9140 7546 9168 7890
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 8956 7398 9076 7426
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 8852 4684 8904 4690
rect 8852 4626 8904 4632
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 8116 4480 8168 4486
rect 8116 4422 8168 4428
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 8760 4480 8812 4486
rect 8760 4422 8812 4428
rect 8128 4146 8156 4422
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 8404 4078 8432 4422
rect 8772 4146 8800 4422
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8576 4072 8628 4078
rect 8864 4026 8892 4626
rect 8576 4014 8628 4020
rect 8220 3836 8516 3856
rect 8276 3834 8300 3836
rect 8356 3834 8380 3836
rect 8436 3834 8460 3836
rect 8298 3782 8300 3834
rect 8362 3782 8374 3834
rect 8436 3782 8438 3834
rect 8276 3780 8300 3782
rect 8356 3780 8380 3782
rect 8436 3780 8460 3782
rect 8220 3760 8516 3780
rect 8300 3664 8352 3670
rect 7668 3624 8300 3652
rect 7104 3596 7156 3602
rect 7104 3538 7156 3544
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 7564 3596 7616 3602
rect 7564 3538 7616 3544
rect 7484 3194 7512 3538
rect 7576 3194 7604 3538
rect 7668 3534 7696 3624
rect 8300 3606 8352 3612
rect 8588 3602 8616 4014
rect 8772 4010 8892 4026
rect 8760 4004 8892 4010
rect 8812 3998 8892 4004
rect 8760 3946 8812 3952
rect 8392 3596 8444 3602
rect 8392 3538 8444 3544
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 8404 3466 8432 3538
rect 8772 3534 8800 3946
rect 8760 3528 8812 3534
rect 8956 3482 8984 7398
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 9048 6662 9076 7278
rect 9416 6798 9444 8298
rect 9508 7478 9536 8366
rect 9692 8090 9720 8463
rect 9784 8294 9812 9472
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 9876 8838 9904 9318
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9772 8288 9824 8294
rect 9772 8230 9824 8236
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9128 6724 9180 6730
rect 9128 6666 9180 6672
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 9048 6186 9076 6598
rect 9140 6361 9168 6666
rect 9508 6662 9536 7414
rect 9968 7410 9996 10406
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 10152 8566 10180 10202
rect 10244 10198 10272 10610
rect 10232 10192 10284 10198
rect 10232 10134 10284 10140
rect 10140 8560 10192 8566
rect 10140 8502 10192 8508
rect 10048 8424 10100 8430
rect 10048 8366 10100 8372
rect 10060 7954 10088 8366
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 10232 8356 10284 8362
rect 10232 8298 10284 8304
rect 10152 8090 10180 8298
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 10244 8022 10272 8298
rect 10232 8016 10284 8022
rect 10232 7958 10284 7964
rect 10048 7948 10100 7954
rect 10048 7890 10100 7896
rect 9956 7404 10008 7410
rect 9956 7346 10008 7352
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9126 6352 9182 6361
rect 9126 6287 9182 6296
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 9036 6180 9088 6186
rect 9036 6122 9088 6128
rect 9048 5846 9076 6122
rect 9036 5840 9088 5846
rect 9036 5782 9088 5788
rect 9034 5672 9090 5681
rect 9034 5607 9036 5616
rect 9088 5607 9090 5616
rect 9036 5578 9088 5584
rect 9140 4758 9168 6190
rect 9588 5568 9640 5574
rect 9586 5536 9588 5545
rect 9640 5536 9642 5545
rect 9586 5471 9642 5480
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 9128 4752 9180 4758
rect 9128 4694 9180 4700
rect 9416 4078 9444 5170
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 8760 3470 8812 3476
rect 8392 3460 8444 3466
rect 8392 3402 8444 3408
rect 8864 3454 8984 3482
rect 8404 3194 8432 3402
rect 8864 3346 8892 3454
rect 8680 3318 8892 3346
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 7564 3188 7616 3194
rect 7564 3130 7616 3136
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 7668 2650 7696 2926
rect 8576 2916 8628 2922
rect 8576 2858 8628 2864
rect 8220 2748 8516 2768
rect 8276 2746 8300 2748
rect 8356 2746 8380 2748
rect 8436 2746 8460 2748
rect 8298 2694 8300 2746
rect 8362 2694 8374 2746
rect 8436 2694 8438 2746
rect 8276 2692 8300 2694
rect 8356 2692 8380 2694
rect 8436 2692 8460 2694
rect 8220 2672 8516 2692
rect 7656 2644 7708 2650
rect 7656 2586 7708 2592
rect 8116 2508 8168 2514
rect 8116 2450 8168 2456
rect 7564 2304 7616 2310
rect 7564 2246 7616 2252
rect 7576 1494 7604 2246
rect 8128 1970 8156 2450
rect 8588 1970 8616 2858
rect 8116 1964 8168 1970
rect 8116 1906 8168 1912
rect 8576 1964 8628 1970
rect 8576 1906 8628 1912
rect 8220 1660 8516 1680
rect 8276 1658 8300 1660
rect 8356 1658 8380 1660
rect 8436 1658 8460 1660
rect 8298 1606 8300 1658
rect 8362 1606 8374 1658
rect 8436 1606 8438 1658
rect 8276 1604 8300 1606
rect 8356 1604 8380 1606
rect 8436 1604 8460 1606
rect 8220 1584 8516 1604
rect 7564 1488 7616 1494
rect 8680 1442 8708 3318
rect 8956 2990 8984 3334
rect 9140 2990 9168 3674
rect 9508 3534 9536 4558
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9324 3126 9352 3334
rect 9312 3120 9364 3126
rect 9312 3062 9364 3068
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 9128 2984 9180 2990
rect 9128 2926 9180 2932
rect 8864 2514 8892 2926
rect 8956 2582 8984 2926
rect 8944 2576 8996 2582
rect 8944 2518 8996 2524
rect 8852 2508 8904 2514
rect 8852 2450 8904 2456
rect 9220 2508 9272 2514
rect 9220 2450 9272 2456
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 8772 1884 8800 2382
rect 9232 2106 9260 2450
rect 9416 2446 9444 2994
rect 9404 2440 9456 2446
rect 9404 2382 9456 2388
rect 9220 2100 9272 2106
rect 9220 2042 9272 2048
rect 8944 1896 8996 1902
rect 8772 1856 8944 1884
rect 8772 1562 8800 1856
rect 8944 1838 8996 1844
rect 8760 1556 8812 1562
rect 8760 1498 8812 1504
rect 7564 1430 7616 1436
rect 8312 1414 8708 1442
rect 9402 1456 9458 1465
rect 8312 800 8340 1414
rect 9402 1391 9404 1400
rect 9456 1391 9458 1400
rect 9404 1362 9456 1368
rect 9692 800 9720 7142
rect 9784 5846 9812 7278
rect 9864 7268 9916 7274
rect 9864 7210 9916 7216
rect 9876 6254 9904 7210
rect 10060 7206 10088 7890
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 10048 7200 10100 7206
rect 10048 7142 10100 7148
rect 9968 6390 9996 7142
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 9956 6384 10008 6390
rect 9956 6326 10008 6332
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9956 6112 10008 6118
rect 9956 6054 10008 6060
rect 9772 5840 9824 5846
rect 9772 5782 9824 5788
rect 9876 5778 9904 6054
rect 9864 5772 9916 5778
rect 9864 5714 9916 5720
rect 9772 5704 9824 5710
rect 9968 5658 9996 6054
rect 9772 5646 9824 5652
rect 9784 5234 9812 5646
rect 9876 5642 9996 5658
rect 9864 5636 9996 5642
rect 9916 5630 9996 5636
rect 9864 5578 9916 5584
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 9864 4684 9916 4690
rect 9864 4626 9916 4632
rect 9772 4548 9824 4554
rect 9772 4490 9824 4496
rect 9784 4146 9812 4490
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9876 3194 9904 4626
rect 10060 4554 10088 6598
rect 10244 5710 10272 7822
rect 10336 7562 10364 12378
rect 10428 12170 10456 12786
rect 10600 12300 10652 12306
rect 10600 12242 10652 12248
rect 10416 12164 10468 12170
rect 10416 12106 10468 12112
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10520 11354 10548 11698
rect 10508 11348 10560 11354
rect 10508 11290 10560 11296
rect 10612 11150 10640 12242
rect 10784 11212 10836 11218
rect 10784 11154 10836 11160
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10416 11008 10468 11014
rect 10416 10950 10468 10956
rect 10600 11008 10652 11014
rect 10600 10950 10652 10956
rect 10428 10470 10456 10950
rect 10612 10674 10640 10950
rect 10508 10668 10560 10674
rect 10508 10610 10560 10616
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10428 9722 10456 10406
rect 10416 9716 10468 9722
rect 10416 9658 10468 9664
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10428 9110 10456 9318
rect 10416 9104 10468 9110
rect 10414 9072 10416 9081
rect 10468 9072 10470 9081
rect 10520 9058 10548 10610
rect 10600 10192 10652 10198
rect 10600 10134 10652 10140
rect 10612 9602 10640 10134
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 10704 9722 10732 9998
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10612 9574 10732 9602
rect 10796 9586 10824 11154
rect 10520 9042 10640 9058
rect 10520 9036 10652 9042
rect 10520 9030 10600 9036
rect 10414 9007 10470 9016
rect 10600 8978 10652 8984
rect 10704 8922 10732 9574
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10796 9178 10824 9318
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 10888 8922 10916 12854
rect 10980 11694 11008 13126
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 10980 11393 11008 11630
rect 10966 11384 11022 11393
rect 10966 11319 11022 11328
rect 10968 11280 11020 11286
rect 10968 11222 11020 11228
rect 10980 10674 11008 11222
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 10980 9353 11008 9454
rect 10966 9344 11022 9353
rect 10966 9279 11022 9288
rect 10612 8894 10732 8922
rect 10796 8894 10916 8922
rect 10508 8560 10560 8566
rect 10508 8502 10560 8508
rect 10416 8288 10468 8294
rect 10416 8230 10468 8236
rect 10428 8090 10456 8230
rect 10416 8084 10468 8090
rect 10416 8026 10468 8032
rect 10520 8022 10548 8502
rect 10508 8016 10560 8022
rect 10508 7958 10560 7964
rect 10612 7886 10640 8894
rect 10690 8528 10746 8537
rect 10690 8463 10692 8472
rect 10744 8463 10746 8472
rect 10692 8434 10744 8440
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10336 7534 10456 7562
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10244 5370 10272 5646
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 10048 4548 10100 4554
rect 10048 4490 10100 4496
rect 10152 3738 10180 4558
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9956 2984 10008 2990
rect 9956 2926 10008 2932
rect 10324 2984 10376 2990
rect 10324 2926 10376 2932
rect 9968 2774 9996 2926
rect 10232 2848 10284 2854
rect 10232 2790 10284 2796
rect 9968 2746 10088 2774
rect 10060 2038 10088 2746
rect 10048 2032 10100 2038
rect 10048 1974 10100 1980
rect 10060 1766 10088 1974
rect 10244 1902 10272 2790
rect 10336 2514 10364 2926
rect 10324 2508 10376 2514
rect 10324 2450 10376 2456
rect 10336 2106 10364 2450
rect 10324 2100 10376 2106
rect 10324 2042 10376 2048
rect 10232 1896 10284 1902
rect 10232 1838 10284 1844
rect 9772 1760 9824 1766
rect 9772 1702 9824 1708
rect 10048 1760 10100 1766
rect 10048 1702 10100 1708
rect 9784 1562 9812 1702
rect 9772 1556 9824 1562
rect 9772 1498 9824 1504
rect 10428 1465 10456 7534
rect 10796 7410 10824 8894
rect 10876 8424 10928 8430
rect 10980 8412 11008 9279
rect 10928 8384 11008 8412
rect 10876 8366 10928 8372
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10888 7546 10916 7686
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10796 6866 10824 7346
rect 10784 6860 10836 6866
rect 10784 6802 10836 6808
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 10508 6656 10560 6662
rect 10508 6598 10560 6604
rect 10520 6254 10548 6598
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10692 6180 10744 6186
rect 10692 6122 10744 6128
rect 10784 6180 10836 6186
rect 10784 6122 10836 6128
rect 10704 5846 10732 6122
rect 10796 5914 10824 6122
rect 10980 5914 11008 6734
rect 10784 5908 10836 5914
rect 10784 5850 10836 5856
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 10692 5840 10744 5846
rect 10692 5782 10744 5788
rect 10796 5370 10824 5850
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 11072 4690 11100 16200
rect 12452 15450 12480 16200
rect 12452 15422 12572 15450
rect 12220 15260 12516 15280
rect 12276 15258 12300 15260
rect 12356 15258 12380 15260
rect 12436 15258 12460 15260
rect 12298 15206 12300 15258
rect 12362 15206 12374 15258
rect 12436 15206 12438 15258
rect 12276 15204 12300 15206
rect 12356 15204 12380 15206
rect 12436 15204 12460 15206
rect 12220 15184 12516 15204
rect 12544 14958 12572 15422
rect 12532 14952 12584 14958
rect 12532 14894 12584 14900
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 11164 10810 11192 14758
rect 12220 14172 12516 14192
rect 12276 14170 12300 14172
rect 12356 14170 12380 14172
rect 12436 14170 12460 14172
rect 12298 14118 12300 14170
rect 12362 14118 12374 14170
rect 12436 14118 12438 14170
rect 12276 14116 12300 14118
rect 12356 14116 12380 14118
rect 12436 14116 12460 14118
rect 12220 14096 12516 14116
rect 11704 14000 11756 14006
rect 11704 13942 11756 13948
rect 11244 13728 11296 13734
rect 11244 13670 11296 13676
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 11256 12850 11284 13670
rect 11624 13394 11652 13670
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 11336 13252 11388 13258
rect 11336 13194 11388 13200
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 11348 12306 11376 13194
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 11164 10606 11192 10746
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 11440 10538 11468 12378
rect 11624 12306 11652 13330
rect 11716 12374 11744 13942
rect 12716 13932 12768 13938
rect 12716 13874 12768 13880
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 11888 13796 11940 13802
rect 11888 13738 11940 13744
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 11704 12368 11756 12374
rect 11704 12310 11756 12316
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11808 11898 11836 12718
rect 11900 12714 11928 13738
rect 12452 13462 12480 13806
rect 12440 13456 12492 13462
rect 12440 13398 12492 13404
rect 12728 13394 12756 13874
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 12992 13728 13044 13734
rect 12992 13670 13044 13676
rect 12716 13388 12768 13394
rect 12716 13330 12768 13336
rect 12220 13084 12516 13104
rect 12276 13082 12300 13084
rect 12356 13082 12380 13084
rect 12436 13082 12460 13084
rect 12298 13030 12300 13082
rect 12362 13030 12374 13082
rect 12436 13030 12438 13082
rect 12276 13028 12300 13030
rect 12356 13028 12380 13030
rect 12436 13028 12460 13030
rect 12220 13008 12516 13028
rect 11888 12708 11940 12714
rect 11888 12650 11940 12656
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11992 11694 12020 12038
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11980 11688 12032 11694
rect 11980 11630 12032 11636
rect 11808 10606 11836 11630
rect 11888 11552 11940 11558
rect 11888 11494 11940 11500
rect 11796 10600 11848 10606
rect 11716 10560 11796 10588
rect 11428 10532 11480 10538
rect 11428 10474 11480 10480
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 11164 9450 11192 10406
rect 11716 10266 11744 10560
rect 11796 10542 11848 10548
rect 11704 10260 11756 10266
rect 11704 10202 11756 10208
rect 11152 9444 11204 9450
rect 11152 9386 11204 9392
rect 11794 9072 11850 9081
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 11336 9036 11388 9042
rect 11794 9007 11796 9016
rect 11336 8978 11388 8984
rect 11848 9007 11850 9016
rect 11796 8978 11848 8984
rect 11164 8906 11192 8978
rect 11152 8900 11204 8906
rect 11152 8842 11204 8848
rect 11348 8634 11376 8978
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 11796 8560 11848 8566
rect 11796 8502 11848 8508
rect 11808 8022 11836 8502
rect 11796 8016 11848 8022
rect 11796 7958 11848 7964
rect 11244 7268 11296 7274
rect 11244 7210 11296 7216
rect 11256 6934 11284 7210
rect 11244 6928 11296 6934
rect 11244 6870 11296 6876
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 11164 5098 11192 6054
rect 11256 5846 11284 6870
rect 11428 6724 11480 6730
rect 11428 6666 11480 6672
rect 11520 6724 11572 6730
rect 11520 6666 11572 6672
rect 11244 5840 11296 5846
rect 11244 5782 11296 5788
rect 11152 5092 11204 5098
rect 11152 5034 11204 5040
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 11060 4684 11112 4690
rect 11060 4626 11112 4632
rect 10612 3602 10640 4626
rect 10692 4616 10744 4622
rect 11072 4570 11100 4626
rect 10692 4558 10744 4564
rect 10704 3602 10732 4558
rect 10980 4542 11100 4570
rect 10980 3602 11008 4542
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 11072 3738 11100 4422
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 10600 3596 10652 3602
rect 10600 3538 10652 3544
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 10612 3505 10640 3538
rect 10598 3496 10654 3505
rect 10598 3431 10654 3440
rect 10612 2496 10640 3431
rect 10704 2650 10732 3538
rect 11060 3188 11112 3194
rect 11060 3130 11112 3136
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 10692 2508 10744 2514
rect 10612 2468 10692 2496
rect 10692 2450 10744 2456
rect 11072 2378 11100 3130
rect 11164 2582 11192 3538
rect 11256 3058 11284 4082
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 11244 2848 11296 2854
rect 11296 2808 11376 2836
rect 11244 2790 11296 2796
rect 11152 2576 11204 2582
rect 11152 2518 11204 2524
rect 11060 2372 11112 2378
rect 11060 2314 11112 2320
rect 11072 2038 11100 2314
rect 11060 2032 11112 2038
rect 11060 1974 11112 1980
rect 11072 1850 11100 1974
rect 11348 1902 11376 2808
rect 10980 1834 11100 1850
rect 11336 1896 11388 1902
rect 11336 1838 11388 1844
rect 10968 1828 11100 1834
rect 11020 1822 11100 1828
rect 10968 1770 11020 1776
rect 10414 1456 10470 1465
rect 11440 1442 11468 6666
rect 11532 5574 11560 6666
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11716 5846 11744 6598
rect 11704 5840 11756 5846
rect 11704 5782 11756 5788
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 11532 4690 11560 5510
rect 11900 5250 11928 11494
rect 11992 11218 12020 11630
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 12084 11121 12112 12174
rect 12808 12164 12860 12170
rect 12808 12106 12860 12112
rect 12220 11996 12516 12016
rect 12276 11994 12300 11996
rect 12356 11994 12380 11996
rect 12436 11994 12460 11996
rect 12298 11942 12300 11994
rect 12362 11942 12374 11994
rect 12436 11942 12438 11994
rect 12276 11940 12300 11942
rect 12356 11940 12380 11942
rect 12436 11940 12460 11942
rect 12220 11920 12516 11940
rect 12820 11762 12848 12106
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 12070 11112 12126 11121
rect 12070 11047 12126 11056
rect 12220 10908 12516 10928
rect 12276 10906 12300 10908
rect 12356 10906 12380 10908
rect 12436 10906 12460 10908
rect 12298 10854 12300 10906
rect 12362 10854 12374 10906
rect 12436 10854 12438 10906
rect 12276 10852 12300 10854
rect 12356 10852 12380 10854
rect 12436 10852 12460 10854
rect 12220 10832 12516 10852
rect 12624 10736 12676 10742
rect 12624 10678 12676 10684
rect 12348 10600 12400 10606
rect 12348 10542 12400 10548
rect 12360 10062 12388 10542
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12072 10056 12124 10062
rect 12072 9998 12124 10004
rect 12348 10056 12400 10062
rect 12348 9998 12400 10004
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11992 9518 12020 9862
rect 12084 9722 12112 9998
rect 12220 9820 12516 9840
rect 12276 9818 12300 9820
rect 12356 9818 12380 9820
rect 12436 9818 12460 9820
rect 12298 9766 12300 9818
rect 12362 9766 12374 9818
rect 12436 9766 12438 9818
rect 12276 9764 12300 9766
rect 12356 9764 12380 9766
rect 12436 9764 12460 9766
rect 12220 9744 12516 9764
rect 12072 9716 12124 9722
rect 12072 9658 12124 9664
rect 11980 9512 12032 9518
rect 11980 9454 12032 9460
rect 11980 8900 12032 8906
rect 11980 8842 12032 8848
rect 11992 6916 12020 8842
rect 12220 8732 12516 8752
rect 12276 8730 12300 8732
rect 12356 8730 12380 8732
rect 12436 8730 12460 8732
rect 12298 8678 12300 8730
rect 12362 8678 12374 8730
rect 12436 8678 12438 8730
rect 12276 8676 12300 8678
rect 12356 8676 12380 8678
rect 12436 8676 12460 8678
rect 12220 8656 12516 8676
rect 12544 8430 12572 10406
rect 12636 9518 12664 10678
rect 12716 10192 12768 10198
rect 12716 10134 12768 10140
rect 12624 9512 12676 9518
rect 12624 9454 12676 9460
rect 12728 9178 12756 10134
rect 12820 9586 12848 11698
rect 13004 10606 13032 13670
rect 13176 13456 13228 13462
rect 13176 13398 13228 13404
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 12992 10600 13044 10606
rect 12992 10542 13044 10548
rect 13004 10130 13032 10542
rect 13096 10198 13124 13126
rect 13188 12782 13216 13398
rect 13176 12776 13228 12782
rect 13176 12718 13228 12724
rect 13188 12442 13216 12718
rect 13176 12436 13228 12442
rect 13176 12378 13228 12384
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 13188 11830 13216 12242
rect 13176 11824 13228 11830
rect 13176 11766 13228 11772
rect 13188 11286 13216 11766
rect 13280 11762 13308 13806
rect 13360 13388 13412 13394
rect 13360 13330 13412 13336
rect 13268 11756 13320 11762
rect 13268 11698 13320 11704
rect 13372 11370 13400 13330
rect 13280 11342 13400 11370
rect 13176 11280 13228 11286
rect 13176 11222 13228 11228
rect 13280 11218 13308 11342
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 13280 10606 13308 11154
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13084 10192 13136 10198
rect 13084 10134 13136 10140
rect 12992 10124 13044 10130
rect 12992 10066 13044 10072
rect 13832 9625 13860 16200
rect 13818 9616 13874 9625
rect 12808 9580 12860 9586
rect 13818 9551 13874 9560
rect 12808 9522 12860 9528
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 12622 8936 12678 8945
rect 12622 8871 12678 8880
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 12636 8362 12664 8871
rect 12820 8498 12848 9522
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 12900 9036 12952 9042
rect 12900 8978 12952 8984
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 12912 8430 12940 8978
rect 12900 8424 12952 8430
rect 12900 8366 12952 8372
rect 12624 8356 12676 8362
rect 12624 8298 12676 8304
rect 12072 8288 12124 8294
rect 12072 8230 12124 8236
rect 12084 7954 12112 8230
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 12084 7342 12112 7890
rect 12220 7644 12516 7664
rect 12276 7642 12300 7644
rect 12356 7642 12380 7644
rect 12436 7642 12460 7644
rect 12298 7590 12300 7642
rect 12362 7590 12374 7642
rect 12436 7590 12438 7642
rect 12276 7588 12300 7590
rect 12356 7588 12380 7590
rect 12436 7588 12460 7590
rect 12220 7568 12516 7588
rect 12072 7336 12124 7342
rect 12072 7278 12124 7284
rect 12440 7336 12492 7342
rect 12492 7284 12572 7290
rect 12440 7278 12572 7284
rect 12452 7262 12572 7278
rect 12072 6928 12124 6934
rect 11992 6888 12072 6916
rect 12072 6870 12124 6876
rect 12220 6556 12516 6576
rect 12276 6554 12300 6556
rect 12356 6554 12380 6556
rect 12436 6554 12460 6556
rect 12298 6502 12300 6554
rect 12362 6502 12374 6554
rect 12436 6502 12438 6554
rect 12276 6500 12300 6502
rect 12356 6500 12380 6502
rect 12436 6500 12460 6502
rect 12220 6480 12516 6500
rect 12220 5468 12516 5488
rect 12276 5466 12300 5468
rect 12356 5466 12380 5468
rect 12436 5466 12460 5468
rect 12298 5414 12300 5466
rect 12362 5414 12374 5466
rect 12436 5414 12438 5466
rect 12276 5412 12300 5414
rect 12356 5412 12380 5414
rect 12436 5412 12460 5414
rect 12220 5392 12516 5412
rect 11900 5222 12020 5250
rect 11888 5160 11940 5166
rect 11888 5102 11940 5108
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 11532 3534 11560 4626
rect 11808 4078 11836 4966
rect 11900 4214 11928 5102
rect 11992 4865 12020 5222
rect 12440 5228 12492 5234
rect 12440 5170 12492 5176
rect 11978 4856 12034 4865
rect 11978 4791 12034 4800
rect 12452 4622 12480 5170
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 12220 4380 12516 4400
rect 12276 4378 12300 4380
rect 12356 4378 12380 4380
rect 12436 4378 12460 4380
rect 12298 4326 12300 4378
rect 12362 4326 12374 4378
rect 12436 4326 12438 4378
rect 12276 4324 12300 4326
rect 12356 4324 12380 4326
rect 12436 4324 12460 4326
rect 12220 4304 12516 4324
rect 11888 4208 11940 4214
rect 11888 4150 11940 4156
rect 11796 4072 11848 4078
rect 11796 4014 11848 4020
rect 11808 3618 11836 4014
rect 11716 3590 11836 3618
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 11532 2582 11560 3470
rect 11716 3058 11744 3590
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 11808 3194 11836 3470
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11900 2990 11928 4150
rect 12072 4004 12124 4010
rect 12072 3946 12124 3952
rect 12084 3482 12112 3946
rect 12544 3618 12572 7262
rect 12716 6792 12768 6798
rect 12716 6734 12768 6740
rect 12728 6322 12756 6734
rect 12716 6316 12768 6322
rect 12716 6258 12768 6264
rect 12912 6254 12940 8366
rect 13360 8016 13412 8022
rect 13360 7958 13412 7964
rect 13268 7948 13320 7954
rect 13268 7890 13320 7896
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 12900 6248 12952 6254
rect 12900 6190 12952 6196
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12820 4758 12848 6054
rect 12808 4752 12860 4758
rect 12808 4694 12860 4700
rect 12912 4214 12940 6190
rect 12900 4208 12952 4214
rect 12900 4150 12952 4156
rect 12900 4072 12952 4078
rect 12900 4014 12952 4020
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12728 3738 12756 3878
rect 12716 3732 12768 3738
rect 12716 3674 12768 3680
rect 12808 3664 12860 3670
rect 12544 3590 12756 3618
rect 12808 3606 12860 3612
rect 12164 3528 12216 3534
rect 12084 3476 12164 3482
rect 12084 3470 12216 3476
rect 12084 3454 12204 3470
rect 11888 2984 11940 2990
rect 11888 2926 11940 2932
rect 11520 2576 11572 2582
rect 11520 2518 11572 2524
rect 10414 1391 10470 1400
rect 11072 1414 11468 1442
rect 11532 1426 11560 2518
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 11624 2106 11652 2382
rect 11796 2304 11848 2310
rect 11900 2258 11928 2926
rect 12084 2922 12112 3454
rect 12220 3292 12516 3312
rect 12276 3290 12300 3292
rect 12356 3290 12380 3292
rect 12436 3290 12460 3292
rect 12298 3238 12300 3290
rect 12362 3238 12374 3290
rect 12436 3238 12438 3290
rect 12276 3236 12300 3238
rect 12356 3236 12380 3238
rect 12436 3236 12460 3238
rect 12220 3216 12516 3236
rect 12532 3120 12584 3126
rect 12532 3062 12584 3068
rect 12072 2916 12124 2922
rect 12072 2858 12124 2864
rect 12256 2848 12308 2854
rect 12256 2790 12308 2796
rect 12268 2650 12296 2790
rect 12256 2644 12308 2650
rect 12256 2586 12308 2592
rect 11848 2252 11928 2258
rect 11796 2246 11928 2252
rect 11808 2230 11928 2246
rect 11612 2100 11664 2106
rect 11612 2042 11664 2048
rect 11900 2038 11928 2230
rect 12220 2204 12516 2224
rect 12276 2202 12300 2204
rect 12356 2202 12380 2204
rect 12436 2202 12460 2204
rect 12298 2150 12300 2202
rect 12362 2150 12374 2202
rect 12436 2150 12438 2202
rect 12276 2148 12300 2150
rect 12356 2148 12380 2150
rect 12436 2148 12460 2150
rect 12220 2128 12516 2148
rect 11888 2032 11940 2038
rect 11888 1974 11940 1980
rect 12256 2032 12308 2038
rect 12256 1974 12308 1980
rect 11520 1420 11572 1426
rect 11072 800 11100 1414
rect 11520 1362 11572 1368
rect 12268 1358 12296 1974
rect 12256 1352 12308 1358
rect 12256 1294 12308 1300
rect 12220 1116 12516 1136
rect 12276 1114 12300 1116
rect 12356 1114 12380 1116
rect 12436 1114 12460 1116
rect 12298 1062 12300 1114
rect 12362 1062 12374 1114
rect 12436 1062 12438 1114
rect 12276 1060 12300 1062
rect 12356 1060 12380 1062
rect 12436 1060 12460 1062
rect 12220 1040 12516 1060
rect 12544 898 12572 3062
rect 12624 2576 12676 2582
rect 12624 2518 12676 2524
rect 12636 1562 12664 2518
rect 12728 2106 12756 3590
rect 12820 3194 12848 3606
rect 12912 3398 12940 4014
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 13004 3194 13032 7346
rect 13082 6896 13138 6905
rect 13082 6831 13138 6840
rect 13096 6798 13124 6831
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 13280 6322 13308 7890
rect 13372 7478 13400 7958
rect 13360 7472 13412 7478
rect 13360 7414 13412 7420
rect 13268 6316 13320 6322
rect 13268 6258 13320 6264
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 13188 5846 13216 6054
rect 13176 5840 13228 5846
rect 13176 5782 13228 5788
rect 13176 5568 13228 5574
rect 13176 5510 13228 5516
rect 13188 5234 13216 5510
rect 13176 5228 13228 5234
rect 13176 5170 13228 5176
rect 13084 5092 13136 5098
rect 13084 5034 13136 5040
rect 13096 4826 13124 5034
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 13084 4072 13136 4078
rect 13084 4014 13136 4020
rect 12808 3188 12860 3194
rect 12808 3130 12860 3136
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 13096 2990 13124 4014
rect 13280 2990 13308 6258
rect 12808 2984 12860 2990
rect 12808 2926 12860 2932
rect 13084 2984 13136 2990
rect 13084 2926 13136 2932
rect 13268 2984 13320 2990
rect 13268 2926 13320 2932
rect 12716 2100 12768 2106
rect 12716 2042 12768 2048
rect 12820 1902 12848 2926
rect 13372 2774 13400 7414
rect 12912 2746 13400 2774
rect 12912 1902 12940 2746
rect 12808 1896 12860 1902
rect 12808 1838 12860 1844
rect 12900 1896 12952 1902
rect 12900 1838 12952 1844
rect 12624 1556 12676 1562
rect 12624 1498 12676 1504
rect 12820 1426 12848 1838
rect 12808 1420 12860 1426
rect 12808 1362 12860 1368
rect 12452 870 12572 898
rect 12452 800 12480 870
rect 13832 800 13860 9318
rect 478 0 534 800
rect 1398 0 1454 800
rect 2778 0 2834 800
rect 4158 0 4214 800
rect 5538 0 5594 800
rect 6918 0 6974 800
rect 8298 0 8354 800
rect 9678 0 9734 800
rect 11058 0 11114 800
rect 12438 0 12494 800
rect 13818 0 13874 800
<< via2 >>
rect 1674 12280 1730 12336
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 4066 14320 4122 14376
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 1858 8200 1914 8256
rect 1858 6160 1914 6216
rect 1858 2080 1914 2136
rect 2686 1420 2742 1456
rect 2686 1400 2688 1420
rect 2688 1400 2740 1420
rect 2740 1400 2742 1420
rect 2870 5652 2872 5672
rect 2872 5652 2924 5672
rect 2924 5652 2926 5672
rect 2870 5616 2926 5652
rect 3514 9560 3570 9616
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 4894 12416 4950 12472
rect 3974 10240 4030 10296
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 3238 4120 3294 4176
rect 5814 12416 5870 12472
rect 5262 6316 5318 6352
rect 5262 6296 5264 6316
rect 5264 6296 5316 6316
rect 5316 6296 5318 6316
rect 8220 15802 8276 15804
rect 8300 15802 8356 15804
rect 8380 15802 8436 15804
rect 8460 15802 8516 15804
rect 8220 15750 8246 15802
rect 8246 15750 8276 15802
rect 8300 15750 8310 15802
rect 8310 15750 8356 15802
rect 8380 15750 8426 15802
rect 8426 15750 8436 15802
rect 8460 15750 8490 15802
rect 8490 15750 8516 15802
rect 8220 15748 8276 15750
rect 8300 15748 8356 15750
rect 8380 15748 8436 15750
rect 8460 15748 8516 15750
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 4220 1114 4276 1116
rect 4300 1114 4356 1116
rect 4380 1114 4436 1116
rect 4460 1114 4516 1116
rect 4220 1062 4246 1114
rect 4246 1062 4276 1114
rect 4300 1062 4310 1114
rect 4310 1062 4356 1114
rect 4380 1062 4426 1114
rect 4426 1062 4436 1114
rect 4460 1062 4490 1114
rect 4490 1062 4516 1114
rect 4220 1060 4276 1062
rect 4300 1060 4356 1062
rect 4380 1060 4436 1062
rect 4460 1060 4516 1062
rect 6550 10124 6606 10160
rect 6550 10104 6552 10124
rect 6552 10104 6604 10124
rect 6604 10104 6606 10124
rect 9862 15020 9918 15056
rect 9862 15000 9864 15020
rect 9864 15000 9916 15020
rect 9916 15000 9918 15020
rect 8220 14714 8276 14716
rect 8300 14714 8356 14716
rect 8380 14714 8436 14716
rect 8460 14714 8516 14716
rect 8220 14662 8246 14714
rect 8246 14662 8276 14714
rect 8300 14662 8310 14714
rect 8310 14662 8356 14714
rect 8380 14662 8426 14714
rect 8426 14662 8436 14714
rect 8460 14662 8490 14714
rect 8490 14662 8516 14714
rect 8220 14660 8276 14662
rect 8300 14660 8356 14662
rect 8380 14660 8436 14662
rect 8460 14660 8516 14662
rect 8220 13626 8276 13628
rect 8300 13626 8356 13628
rect 8380 13626 8436 13628
rect 8460 13626 8516 13628
rect 8220 13574 8246 13626
rect 8246 13574 8276 13626
rect 8300 13574 8310 13626
rect 8310 13574 8356 13626
rect 8380 13574 8426 13626
rect 8426 13574 8436 13626
rect 8460 13574 8490 13626
rect 8490 13574 8516 13626
rect 8220 13572 8276 13574
rect 8300 13572 8356 13574
rect 8380 13572 8436 13574
rect 8460 13572 8516 13574
rect 8220 12538 8276 12540
rect 8300 12538 8356 12540
rect 8380 12538 8436 12540
rect 8460 12538 8516 12540
rect 8220 12486 8246 12538
rect 8246 12486 8276 12538
rect 8300 12486 8310 12538
rect 8310 12486 8356 12538
rect 8380 12486 8426 12538
rect 8426 12486 8436 12538
rect 8460 12486 8490 12538
rect 8490 12486 8516 12538
rect 8220 12484 8276 12486
rect 8300 12484 8356 12486
rect 8380 12484 8436 12486
rect 8460 12484 8516 12486
rect 8482 12144 8538 12200
rect 8482 11600 8538 11656
rect 8022 10124 8078 10160
rect 8220 11450 8276 11452
rect 8300 11450 8356 11452
rect 8380 11450 8436 11452
rect 8460 11450 8516 11452
rect 8220 11398 8246 11450
rect 8246 11398 8276 11450
rect 8300 11398 8310 11450
rect 8310 11398 8356 11450
rect 8380 11398 8426 11450
rect 8426 11398 8436 11450
rect 8460 11398 8490 11450
rect 8490 11398 8516 11450
rect 8220 11396 8276 11398
rect 8300 11396 8356 11398
rect 8380 11396 8436 11398
rect 8460 11396 8516 11398
rect 8220 10362 8276 10364
rect 8300 10362 8356 10364
rect 8380 10362 8436 10364
rect 8460 10362 8516 10364
rect 8220 10310 8246 10362
rect 8246 10310 8276 10362
rect 8300 10310 8310 10362
rect 8310 10310 8356 10362
rect 8380 10310 8426 10362
rect 8426 10310 8436 10362
rect 8460 10310 8490 10362
rect 8490 10310 8516 10362
rect 8220 10308 8276 10310
rect 8300 10308 8356 10310
rect 8380 10308 8436 10310
rect 8460 10308 8516 10310
rect 8022 10104 8024 10124
rect 8024 10104 8076 10124
rect 8076 10104 8078 10124
rect 8022 9424 8078 9480
rect 7654 7384 7710 7440
rect 8220 9274 8276 9276
rect 8300 9274 8356 9276
rect 8380 9274 8436 9276
rect 8460 9274 8516 9276
rect 8220 9222 8246 9274
rect 8246 9222 8276 9274
rect 8300 9222 8310 9274
rect 8310 9222 8356 9274
rect 8380 9222 8426 9274
rect 8426 9222 8436 9274
rect 8460 9222 8490 9274
rect 8490 9222 8516 9274
rect 8220 9220 8276 9222
rect 8300 9220 8356 9222
rect 8380 9220 8436 9222
rect 8460 9220 8516 9222
rect 8220 8186 8276 8188
rect 8300 8186 8356 8188
rect 8380 8186 8436 8188
rect 8460 8186 8516 8188
rect 8220 8134 8246 8186
rect 8246 8134 8276 8186
rect 8300 8134 8310 8186
rect 8310 8134 8356 8186
rect 8380 8134 8426 8186
rect 8426 8134 8436 8186
rect 8460 8134 8490 8186
rect 8490 8134 8516 8186
rect 8220 8132 8276 8134
rect 8300 8132 8356 8134
rect 8380 8132 8436 8134
rect 8460 8132 8516 8134
rect 8022 7792 8078 7848
rect 8220 7098 8276 7100
rect 8300 7098 8356 7100
rect 8380 7098 8436 7100
rect 8460 7098 8516 7100
rect 8220 7046 8246 7098
rect 8246 7046 8276 7098
rect 8300 7046 8310 7098
rect 8310 7046 8356 7098
rect 8380 7046 8426 7098
rect 8426 7046 8436 7098
rect 8460 7046 8490 7098
rect 8490 7046 8516 7098
rect 8220 7044 8276 7046
rect 8300 7044 8356 7046
rect 8380 7044 8436 7046
rect 8460 7044 8516 7046
rect 8220 6010 8276 6012
rect 8300 6010 8356 6012
rect 8380 6010 8436 6012
rect 8460 6010 8516 6012
rect 8220 5958 8246 6010
rect 8246 5958 8276 6010
rect 8300 5958 8310 6010
rect 8310 5958 8356 6010
rect 8380 5958 8426 6010
rect 8426 5958 8436 6010
rect 8460 5958 8490 6010
rect 8490 5958 8516 6010
rect 8220 5956 8276 5958
rect 8300 5956 8356 5958
rect 8380 5956 8436 5958
rect 8460 5956 8516 5958
rect 8482 5516 8484 5536
rect 8484 5516 8536 5536
rect 8536 5516 8538 5536
rect 8482 5480 8538 5516
rect 8220 4922 8276 4924
rect 8300 4922 8356 4924
rect 8380 4922 8436 4924
rect 8460 4922 8516 4924
rect 8220 4870 8246 4922
rect 8246 4870 8276 4922
rect 8300 4870 8310 4922
rect 8310 4870 8356 4922
rect 8380 4870 8426 4922
rect 8426 4870 8436 4922
rect 8460 4870 8490 4922
rect 8490 4870 8516 4922
rect 8220 4868 8276 4870
rect 8300 4868 8356 4870
rect 8380 4868 8436 4870
rect 8460 4868 8516 4870
rect 9218 11600 9274 11656
rect 9586 11600 9642 11656
rect 9402 11328 9458 11384
rect 9862 12144 9918 12200
rect 9586 9424 9642 9480
rect 9678 9288 9734 9344
rect 9678 8472 9734 8528
rect 8220 3834 8276 3836
rect 8300 3834 8356 3836
rect 8380 3834 8436 3836
rect 8460 3834 8516 3836
rect 8220 3782 8246 3834
rect 8246 3782 8276 3834
rect 8300 3782 8310 3834
rect 8310 3782 8356 3834
rect 8380 3782 8426 3834
rect 8426 3782 8436 3834
rect 8460 3782 8490 3834
rect 8490 3782 8516 3834
rect 8220 3780 8276 3782
rect 8300 3780 8356 3782
rect 8380 3780 8436 3782
rect 8460 3780 8516 3782
rect 9126 6296 9182 6352
rect 9034 5636 9090 5672
rect 9034 5616 9036 5636
rect 9036 5616 9088 5636
rect 9088 5616 9090 5636
rect 9586 5516 9588 5536
rect 9588 5516 9640 5536
rect 9640 5516 9642 5536
rect 9586 5480 9642 5516
rect 8220 2746 8276 2748
rect 8300 2746 8356 2748
rect 8380 2746 8436 2748
rect 8460 2746 8516 2748
rect 8220 2694 8246 2746
rect 8246 2694 8276 2746
rect 8300 2694 8310 2746
rect 8310 2694 8356 2746
rect 8380 2694 8426 2746
rect 8426 2694 8436 2746
rect 8460 2694 8490 2746
rect 8490 2694 8516 2746
rect 8220 2692 8276 2694
rect 8300 2692 8356 2694
rect 8380 2692 8436 2694
rect 8460 2692 8516 2694
rect 8220 1658 8276 1660
rect 8300 1658 8356 1660
rect 8380 1658 8436 1660
rect 8460 1658 8516 1660
rect 8220 1606 8246 1658
rect 8246 1606 8276 1658
rect 8300 1606 8310 1658
rect 8310 1606 8356 1658
rect 8380 1606 8426 1658
rect 8426 1606 8436 1658
rect 8460 1606 8490 1658
rect 8490 1606 8516 1658
rect 8220 1604 8276 1606
rect 8300 1604 8356 1606
rect 8380 1604 8436 1606
rect 8460 1604 8516 1606
rect 9402 1420 9458 1456
rect 9402 1400 9404 1420
rect 9404 1400 9456 1420
rect 9456 1400 9458 1420
rect 10414 9052 10416 9072
rect 10416 9052 10468 9072
rect 10468 9052 10470 9072
rect 10414 9016 10470 9052
rect 10966 11328 11022 11384
rect 10966 9288 11022 9344
rect 10690 8492 10746 8528
rect 10690 8472 10692 8492
rect 10692 8472 10744 8492
rect 10744 8472 10746 8492
rect 12220 15258 12276 15260
rect 12300 15258 12356 15260
rect 12380 15258 12436 15260
rect 12460 15258 12516 15260
rect 12220 15206 12246 15258
rect 12246 15206 12276 15258
rect 12300 15206 12310 15258
rect 12310 15206 12356 15258
rect 12380 15206 12426 15258
rect 12426 15206 12436 15258
rect 12460 15206 12490 15258
rect 12490 15206 12516 15258
rect 12220 15204 12276 15206
rect 12300 15204 12356 15206
rect 12380 15204 12436 15206
rect 12460 15204 12516 15206
rect 12220 14170 12276 14172
rect 12300 14170 12356 14172
rect 12380 14170 12436 14172
rect 12460 14170 12516 14172
rect 12220 14118 12246 14170
rect 12246 14118 12276 14170
rect 12300 14118 12310 14170
rect 12310 14118 12356 14170
rect 12380 14118 12426 14170
rect 12426 14118 12436 14170
rect 12460 14118 12490 14170
rect 12490 14118 12516 14170
rect 12220 14116 12276 14118
rect 12300 14116 12356 14118
rect 12380 14116 12436 14118
rect 12460 14116 12516 14118
rect 12220 13082 12276 13084
rect 12300 13082 12356 13084
rect 12380 13082 12436 13084
rect 12460 13082 12516 13084
rect 12220 13030 12246 13082
rect 12246 13030 12276 13082
rect 12300 13030 12310 13082
rect 12310 13030 12356 13082
rect 12380 13030 12426 13082
rect 12426 13030 12436 13082
rect 12460 13030 12490 13082
rect 12490 13030 12516 13082
rect 12220 13028 12276 13030
rect 12300 13028 12356 13030
rect 12380 13028 12436 13030
rect 12460 13028 12516 13030
rect 11794 9036 11850 9072
rect 11794 9016 11796 9036
rect 11796 9016 11848 9036
rect 11848 9016 11850 9036
rect 10598 3440 10654 3496
rect 10414 1400 10470 1456
rect 12220 11994 12276 11996
rect 12300 11994 12356 11996
rect 12380 11994 12436 11996
rect 12460 11994 12516 11996
rect 12220 11942 12246 11994
rect 12246 11942 12276 11994
rect 12300 11942 12310 11994
rect 12310 11942 12356 11994
rect 12380 11942 12426 11994
rect 12426 11942 12436 11994
rect 12460 11942 12490 11994
rect 12490 11942 12516 11994
rect 12220 11940 12276 11942
rect 12300 11940 12356 11942
rect 12380 11940 12436 11942
rect 12460 11940 12516 11942
rect 12070 11056 12126 11112
rect 12220 10906 12276 10908
rect 12300 10906 12356 10908
rect 12380 10906 12436 10908
rect 12460 10906 12516 10908
rect 12220 10854 12246 10906
rect 12246 10854 12276 10906
rect 12300 10854 12310 10906
rect 12310 10854 12356 10906
rect 12380 10854 12426 10906
rect 12426 10854 12436 10906
rect 12460 10854 12490 10906
rect 12490 10854 12516 10906
rect 12220 10852 12276 10854
rect 12300 10852 12356 10854
rect 12380 10852 12436 10854
rect 12460 10852 12516 10854
rect 12220 9818 12276 9820
rect 12300 9818 12356 9820
rect 12380 9818 12436 9820
rect 12460 9818 12516 9820
rect 12220 9766 12246 9818
rect 12246 9766 12276 9818
rect 12300 9766 12310 9818
rect 12310 9766 12356 9818
rect 12380 9766 12426 9818
rect 12426 9766 12436 9818
rect 12460 9766 12490 9818
rect 12490 9766 12516 9818
rect 12220 9764 12276 9766
rect 12300 9764 12356 9766
rect 12380 9764 12436 9766
rect 12460 9764 12516 9766
rect 12220 8730 12276 8732
rect 12300 8730 12356 8732
rect 12380 8730 12436 8732
rect 12460 8730 12516 8732
rect 12220 8678 12246 8730
rect 12246 8678 12276 8730
rect 12300 8678 12310 8730
rect 12310 8678 12356 8730
rect 12380 8678 12426 8730
rect 12426 8678 12436 8730
rect 12460 8678 12490 8730
rect 12490 8678 12516 8730
rect 12220 8676 12276 8678
rect 12300 8676 12356 8678
rect 12380 8676 12436 8678
rect 12460 8676 12516 8678
rect 13818 9560 13874 9616
rect 12622 8880 12678 8936
rect 12220 7642 12276 7644
rect 12300 7642 12356 7644
rect 12380 7642 12436 7644
rect 12460 7642 12516 7644
rect 12220 7590 12246 7642
rect 12246 7590 12276 7642
rect 12300 7590 12310 7642
rect 12310 7590 12356 7642
rect 12380 7590 12426 7642
rect 12426 7590 12436 7642
rect 12460 7590 12490 7642
rect 12490 7590 12516 7642
rect 12220 7588 12276 7590
rect 12300 7588 12356 7590
rect 12380 7588 12436 7590
rect 12460 7588 12516 7590
rect 12220 6554 12276 6556
rect 12300 6554 12356 6556
rect 12380 6554 12436 6556
rect 12460 6554 12516 6556
rect 12220 6502 12246 6554
rect 12246 6502 12276 6554
rect 12300 6502 12310 6554
rect 12310 6502 12356 6554
rect 12380 6502 12426 6554
rect 12426 6502 12436 6554
rect 12460 6502 12490 6554
rect 12490 6502 12516 6554
rect 12220 6500 12276 6502
rect 12300 6500 12356 6502
rect 12380 6500 12436 6502
rect 12460 6500 12516 6502
rect 12220 5466 12276 5468
rect 12300 5466 12356 5468
rect 12380 5466 12436 5468
rect 12460 5466 12516 5468
rect 12220 5414 12246 5466
rect 12246 5414 12276 5466
rect 12300 5414 12310 5466
rect 12310 5414 12356 5466
rect 12380 5414 12426 5466
rect 12426 5414 12436 5466
rect 12460 5414 12490 5466
rect 12490 5414 12516 5466
rect 12220 5412 12276 5414
rect 12300 5412 12356 5414
rect 12380 5412 12436 5414
rect 12460 5412 12516 5414
rect 11978 4800 12034 4856
rect 12220 4378 12276 4380
rect 12300 4378 12356 4380
rect 12380 4378 12436 4380
rect 12460 4378 12516 4380
rect 12220 4326 12246 4378
rect 12246 4326 12276 4378
rect 12300 4326 12310 4378
rect 12310 4326 12356 4378
rect 12380 4326 12426 4378
rect 12426 4326 12436 4378
rect 12460 4326 12490 4378
rect 12490 4326 12516 4378
rect 12220 4324 12276 4326
rect 12300 4324 12356 4326
rect 12380 4324 12436 4326
rect 12460 4324 12516 4326
rect 12220 3290 12276 3292
rect 12300 3290 12356 3292
rect 12380 3290 12436 3292
rect 12460 3290 12516 3292
rect 12220 3238 12246 3290
rect 12246 3238 12276 3290
rect 12300 3238 12310 3290
rect 12310 3238 12356 3290
rect 12380 3238 12426 3290
rect 12426 3238 12436 3290
rect 12460 3238 12490 3290
rect 12490 3238 12516 3290
rect 12220 3236 12276 3238
rect 12300 3236 12356 3238
rect 12380 3236 12436 3238
rect 12460 3236 12516 3238
rect 12220 2202 12276 2204
rect 12300 2202 12356 2204
rect 12380 2202 12436 2204
rect 12460 2202 12516 2204
rect 12220 2150 12246 2202
rect 12246 2150 12276 2202
rect 12300 2150 12310 2202
rect 12310 2150 12356 2202
rect 12380 2150 12426 2202
rect 12426 2150 12436 2202
rect 12460 2150 12490 2202
rect 12490 2150 12516 2202
rect 12220 2148 12276 2150
rect 12300 2148 12356 2150
rect 12380 2148 12436 2150
rect 12460 2148 12516 2150
rect 12220 1114 12276 1116
rect 12300 1114 12356 1116
rect 12380 1114 12436 1116
rect 12460 1114 12516 1116
rect 12220 1062 12246 1114
rect 12246 1062 12276 1114
rect 12300 1062 12310 1114
rect 12310 1062 12356 1114
rect 12380 1062 12426 1114
rect 12426 1062 12436 1114
rect 12460 1062 12490 1114
rect 12490 1062 12516 1114
rect 12220 1060 12276 1062
rect 12300 1060 12356 1062
rect 12380 1060 12436 1062
rect 12460 1060 12516 1062
rect 13082 6840 13138 6896
<< metal3 >>
rect 8208 15808 8528 15809
rect 8208 15744 8216 15808
rect 8280 15744 8296 15808
rect 8360 15744 8376 15808
rect 8440 15744 8456 15808
rect 8520 15744 8528 15808
rect 8208 15743 8528 15744
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 12208 15264 12528 15265
rect 12208 15200 12216 15264
rect 12280 15200 12296 15264
rect 12360 15200 12376 15264
rect 12440 15200 12456 15264
rect 12520 15200 12528 15264
rect 12208 15199 12528 15200
rect 9857 15058 9923 15061
rect 14200 15058 15000 15088
rect 9857 15056 15000 15058
rect 9857 15000 9862 15056
rect 9918 15000 15000 15056
rect 9857 14998 15000 15000
rect 9857 14995 9923 14998
rect 14200 14968 15000 14998
rect 8208 14720 8528 14721
rect 8208 14656 8216 14720
rect 8280 14656 8296 14720
rect 8360 14656 8376 14720
rect 8440 14656 8456 14720
rect 8520 14656 8528 14720
rect 8208 14655 8528 14656
rect 0 14378 800 14408
rect 4061 14378 4127 14381
rect 0 14376 4127 14378
rect 0 14320 4066 14376
rect 4122 14320 4127 14376
rect 0 14318 4127 14320
rect 0 14288 800 14318
rect 4061 14315 4127 14318
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 12208 14176 12528 14177
rect 12208 14112 12216 14176
rect 12280 14112 12296 14176
rect 12360 14112 12376 14176
rect 12440 14112 12456 14176
rect 12520 14112 12528 14176
rect 12208 14111 12528 14112
rect 8208 13632 8528 13633
rect 8208 13568 8216 13632
rect 8280 13568 8296 13632
rect 8360 13568 8376 13632
rect 8440 13568 8456 13632
rect 8520 13568 8528 13632
rect 8208 13567 8528 13568
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 12208 13088 12528 13089
rect 12208 13024 12216 13088
rect 12280 13024 12296 13088
rect 12360 13024 12376 13088
rect 12440 13024 12456 13088
rect 12520 13024 12528 13088
rect 12208 13023 12528 13024
rect 14200 12928 15000 13048
rect 8208 12544 8528 12545
rect 8208 12480 8216 12544
rect 8280 12480 8296 12544
rect 8360 12480 8376 12544
rect 8440 12480 8456 12544
rect 8520 12480 8528 12544
rect 8208 12479 8528 12480
rect 4889 12474 4955 12477
rect 5809 12474 5875 12477
rect 4889 12472 5875 12474
rect 4889 12416 4894 12472
rect 4950 12416 5814 12472
rect 5870 12416 5875 12472
rect 4889 12414 5875 12416
rect 4889 12411 4955 12414
rect 5809 12411 5875 12414
rect 0 12338 800 12368
rect 1669 12338 1735 12341
rect 0 12336 1735 12338
rect 0 12280 1674 12336
rect 1730 12280 1735 12336
rect 0 12278 1735 12280
rect 0 12248 800 12278
rect 1669 12275 1735 12278
rect 8477 12202 8543 12205
rect 9857 12202 9923 12205
rect 8477 12200 9923 12202
rect 8477 12144 8482 12200
rect 8538 12144 9862 12200
rect 9918 12144 9923 12200
rect 8477 12142 9923 12144
rect 8477 12139 8543 12142
rect 9857 12139 9923 12142
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 12208 12000 12528 12001
rect 12208 11936 12216 12000
rect 12280 11936 12296 12000
rect 12360 11936 12376 12000
rect 12440 11936 12456 12000
rect 12520 11936 12528 12000
rect 12208 11935 12528 11936
rect 8477 11658 8543 11661
rect 9213 11658 9279 11661
rect 9581 11658 9647 11661
rect 8477 11656 9647 11658
rect 8477 11600 8482 11656
rect 8538 11600 9218 11656
rect 9274 11600 9586 11656
rect 9642 11600 9647 11656
rect 8477 11598 9647 11600
rect 8477 11595 8543 11598
rect 9213 11595 9279 11598
rect 9581 11595 9647 11598
rect 8208 11456 8528 11457
rect 8208 11392 8216 11456
rect 8280 11392 8296 11456
rect 8360 11392 8376 11456
rect 8440 11392 8456 11456
rect 8520 11392 8528 11456
rect 8208 11391 8528 11392
rect 9397 11386 9463 11389
rect 10961 11386 11027 11389
rect 9397 11384 11027 11386
rect 9397 11328 9402 11384
rect 9458 11328 10966 11384
rect 11022 11328 11027 11384
rect 9397 11326 11027 11328
rect 9397 11323 9463 11326
rect 10961 11323 11027 11326
rect 12065 11114 12131 11117
rect 12065 11112 12818 11114
rect 12065 11056 12070 11112
rect 12126 11056 12818 11112
rect 12065 11054 12818 11056
rect 12065 11051 12131 11054
rect 12758 10978 12818 11054
rect 14200 10978 15000 11008
rect 12758 10918 15000 10978
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 12208 10912 12528 10913
rect 12208 10848 12216 10912
rect 12280 10848 12296 10912
rect 12360 10848 12376 10912
rect 12440 10848 12456 10912
rect 12520 10848 12528 10912
rect 14200 10888 15000 10918
rect 12208 10847 12528 10848
rect 8208 10368 8528 10369
rect 0 10298 800 10328
rect 8208 10304 8216 10368
rect 8280 10304 8296 10368
rect 8360 10304 8376 10368
rect 8440 10304 8456 10368
rect 8520 10304 8528 10368
rect 8208 10303 8528 10304
rect 3969 10298 4035 10301
rect 0 10296 4035 10298
rect 0 10240 3974 10296
rect 4030 10240 4035 10296
rect 0 10238 4035 10240
rect 0 10208 800 10238
rect 3969 10235 4035 10238
rect 6545 10162 6611 10165
rect 8017 10162 8083 10165
rect 6545 10160 8083 10162
rect 6545 10104 6550 10160
rect 6606 10104 8022 10160
rect 8078 10104 8083 10160
rect 6545 10102 8083 10104
rect 6545 10099 6611 10102
rect 8017 10099 8083 10102
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 12208 9824 12528 9825
rect 12208 9760 12216 9824
rect 12280 9760 12296 9824
rect 12360 9760 12376 9824
rect 12440 9760 12456 9824
rect 12520 9760 12528 9824
rect 12208 9759 12528 9760
rect 3509 9618 3575 9621
rect 13813 9618 13879 9621
rect 3509 9616 13879 9618
rect 3509 9560 3514 9616
rect 3570 9560 13818 9616
rect 13874 9560 13879 9616
rect 3509 9558 13879 9560
rect 3509 9555 3575 9558
rect 13813 9555 13879 9558
rect 8017 9482 8083 9485
rect 9581 9482 9647 9485
rect 8017 9480 9647 9482
rect 8017 9424 8022 9480
rect 8078 9424 9586 9480
rect 9642 9424 9647 9480
rect 8017 9422 9647 9424
rect 8017 9419 8083 9422
rect 9581 9419 9647 9422
rect 9673 9346 9739 9349
rect 10961 9346 11027 9349
rect 9673 9344 11027 9346
rect 9673 9288 9678 9344
rect 9734 9288 10966 9344
rect 11022 9288 11027 9344
rect 9673 9286 11027 9288
rect 9673 9283 9739 9286
rect 10961 9283 11027 9286
rect 8208 9280 8528 9281
rect 8208 9216 8216 9280
rect 8280 9216 8296 9280
rect 8360 9216 8376 9280
rect 8440 9216 8456 9280
rect 8520 9216 8528 9280
rect 8208 9215 8528 9216
rect 10409 9074 10475 9077
rect 11789 9074 11855 9077
rect 10409 9072 11855 9074
rect 10409 9016 10414 9072
rect 10470 9016 11794 9072
rect 11850 9016 11855 9072
rect 10409 9014 11855 9016
rect 10409 9011 10475 9014
rect 11789 9011 11855 9014
rect 12617 8938 12683 8941
rect 14200 8938 15000 8968
rect 12617 8936 15000 8938
rect 12617 8880 12622 8936
rect 12678 8880 15000 8936
rect 12617 8878 15000 8880
rect 12617 8875 12683 8878
rect 14200 8848 15000 8878
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 12208 8736 12528 8737
rect 12208 8672 12216 8736
rect 12280 8672 12296 8736
rect 12360 8672 12376 8736
rect 12440 8672 12456 8736
rect 12520 8672 12528 8736
rect 12208 8671 12528 8672
rect 9673 8530 9739 8533
rect 10685 8530 10751 8533
rect 9673 8528 10751 8530
rect 9673 8472 9678 8528
rect 9734 8472 10690 8528
rect 10746 8472 10751 8528
rect 9673 8470 10751 8472
rect 9673 8467 9739 8470
rect 10685 8467 10751 8470
rect 0 8258 800 8288
rect 1853 8258 1919 8261
rect 0 8256 1919 8258
rect 0 8200 1858 8256
rect 1914 8200 1919 8256
rect 0 8198 1919 8200
rect 0 8168 800 8198
rect 1853 8195 1919 8198
rect 8208 8192 8528 8193
rect 8208 8128 8216 8192
rect 8280 8128 8296 8192
rect 8360 8128 8376 8192
rect 8440 8128 8456 8192
rect 8520 8128 8528 8192
rect 8208 8127 8528 8128
rect 8017 7850 8083 7853
rect 7974 7848 8083 7850
rect 7974 7792 8022 7848
rect 8078 7792 8083 7848
rect 7974 7787 8083 7792
rect 4210 7649 4524 7656
rect 4208 7644 4528 7649
rect 4208 7588 4220 7644
rect 4276 7588 4300 7644
rect 4356 7588 4380 7644
rect 4436 7588 4460 7644
rect 4516 7588 4528 7644
rect 4208 7583 4528 7588
rect 4210 7580 4524 7583
rect 7649 7442 7715 7445
rect 7974 7442 8034 7787
rect 12210 7649 12524 7654
rect 12208 7644 12528 7649
rect 12208 7588 12220 7644
rect 12276 7588 12300 7644
rect 12356 7588 12380 7644
rect 12436 7588 12460 7644
rect 12516 7588 12528 7644
rect 12208 7583 12528 7588
rect 12210 7578 12524 7583
rect 7649 7440 8034 7442
rect 7649 7384 7654 7440
rect 7710 7384 8034 7440
rect 7649 7382 8034 7384
rect 7649 7379 7715 7382
rect 8208 7104 8528 7105
rect 8208 7040 8216 7104
rect 8280 7040 8296 7104
rect 8360 7040 8376 7104
rect 8440 7040 8456 7104
rect 8520 7040 8528 7104
rect 8208 7039 8528 7040
rect 13077 6898 13143 6901
rect 14200 6898 15000 6928
rect 13077 6896 15000 6898
rect 13077 6840 13082 6896
rect 13138 6840 15000 6896
rect 13077 6838 15000 6840
rect 13077 6835 13143 6838
rect 14200 6808 15000 6838
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 12208 6560 12528 6561
rect 12208 6496 12216 6560
rect 12280 6496 12296 6560
rect 12360 6496 12376 6560
rect 12440 6496 12456 6560
rect 12520 6496 12528 6560
rect 12208 6495 12528 6496
rect 5257 6354 5323 6357
rect 9121 6354 9187 6357
rect 5257 6352 9187 6354
rect 5257 6296 5262 6352
rect 5318 6296 9126 6352
rect 9182 6296 9187 6352
rect 5257 6294 9187 6296
rect 5257 6291 5323 6294
rect 9121 6291 9187 6294
rect 0 6218 800 6248
rect 1853 6218 1919 6221
rect 0 6216 1919 6218
rect 0 6160 1858 6216
rect 1914 6160 1919 6216
rect 0 6158 1919 6160
rect 0 6128 800 6158
rect 1853 6155 1919 6158
rect 8208 6016 8528 6017
rect 8208 5952 8216 6016
rect 8280 5952 8296 6016
rect 8360 5952 8376 6016
rect 8440 5952 8456 6016
rect 8520 5952 8528 6016
rect 8208 5951 8528 5952
rect 2865 5674 2931 5677
rect 9029 5674 9095 5677
rect 2865 5672 9095 5674
rect 2865 5616 2870 5672
rect 2926 5616 9034 5672
rect 9090 5616 9095 5672
rect 2865 5614 9095 5616
rect 2865 5611 2931 5614
rect 9029 5611 9095 5614
rect 8477 5538 8543 5541
rect 9581 5538 9647 5541
rect 8477 5536 9647 5538
rect 8477 5480 8482 5536
rect 8538 5480 9586 5536
rect 9642 5480 9647 5536
rect 8477 5478 9647 5480
rect 8477 5475 8543 5478
rect 9581 5475 9647 5478
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 12208 5472 12528 5473
rect 12208 5408 12216 5472
rect 12280 5408 12296 5472
rect 12360 5408 12376 5472
rect 12440 5408 12456 5472
rect 12520 5408 12528 5472
rect 12208 5407 12528 5408
rect 8208 4928 8528 4929
rect 8208 4864 8216 4928
rect 8280 4864 8296 4928
rect 8360 4864 8376 4928
rect 8440 4864 8456 4928
rect 8520 4864 8528 4928
rect 8208 4863 8528 4864
rect 11973 4858 12039 4861
rect 14200 4858 15000 4888
rect 11973 4856 15000 4858
rect 11973 4800 11978 4856
rect 12034 4800 15000 4856
rect 11973 4798 15000 4800
rect 11973 4795 12039 4798
rect 14200 4768 15000 4798
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 12208 4384 12528 4385
rect 12208 4320 12216 4384
rect 12280 4320 12296 4384
rect 12360 4320 12376 4384
rect 12440 4320 12456 4384
rect 12520 4320 12528 4384
rect 12208 4319 12528 4320
rect 0 4178 800 4208
rect 3233 4178 3299 4181
rect 0 4176 3299 4178
rect 0 4120 3238 4176
rect 3294 4120 3299 4176
rect 0 4118 3299 4120
rect 0 4088 800 4118
rect 3233 4115 3299 4118
rect 8208 3840 8528 3841
rect 8208 3776 8216 3840
rect 8280 3776 8296 3840
rect 8360 3776 8376 3840
rect 8440 3776 8456 3840
rect 8520 3776 8528 3840
rect 8208 3775 8528 3776
rect 10593 3498 10659 3501
rect 14200 3498 15000 3528
rect 10593 3496 15000 3498
rect 10593 3440 10598 3496
rect 10654 3440 15000 3496
rect 10593 3438 15000 3440
rect 10593 3435 10659 3438
rect 14200 3408 15000 3438
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 12208 3296 12528 3297
rect 12208 3232 12216 3296
rect 12280 3232 12296 3296
rect 12360 3232 12376 3296
rect 12440 3232 12456 3296
rect 12520 3232 12528 3296
rect 12208 3231 12528 3232
rect 8208 2752 8528 2753
rect 8208 2688 8216 2752
rect 8280 2688 8296 2752
rect 8360 2688 8376 2752
rect 8440 2688 8456 2752
rect 8520 2688 8528 2752
rect 8208 2687 8528 2688
rect 4208 2208 4528 2209
rect 0 2138 800 2168
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 12208 2208 12528 2209
rect 12208 2144 12216 2208
rect 12280 2144 12296 2208
rect 12360 2144 12376 2208
rect 12440 2144 12456 2208
rect 12520 2144 12528 2208
rect 12208 2143 12528 2144
rect 1853 2138 1919 2141
rect 0 2136 1919 2138
rect 0 2080 1858 2136
rect 1914 2080 1919 2136
rect 0 2078 1919 2080
rect 0 2048 800 2078
rect 1853 2075 1919 2078
rect 8208 1664 8528 1665
rect 8208 1600 8216 1664
rect 8280 1600 8296 1664
rect 8360 1600 8376 1664
rect 8440 1600 8456 1664
rect 8520 1600 8528 1664
rect 8208 1599 8528 1600
rect 2681 1458 2747 1461
rect 9397 1458 9463 1461
rect 2681 1456 9463 1458
rect 2681 1400 2686 1456
rect 2742 1400 9402 1456
rect 9458 1400 9463 1456
rect 2681 1398 9463 1400
rect 2681 1395 2747 1398
rect 9397 1395 9463 1398
rect 10409 1458 10475 1461
rect 14200 1458 15000 1488
rect 10409 1456 15000 1458
rect 10409 1400 10414 1456
rect 10470 1400 15000 1456
rect 10409 1398 15000 1400
rect 10409 1395 10475 1398
rect 14200 1368 15000 1398
rect 4208 1120 4528 1121
rect 4208 1056 4216 1120
rect 4280 1056 4296 1120
rect 4360 1056 4376 1120
rect 4440 1056 4456 1120
rect 4520 1056 4528 1120
rect 4208 1055 4528 1056
rect 12208 1120 12528 1121
rect 12208 1056 12216 1120
rect 12280 1056 12296 1120
rect 12360 1056 12376 1120
rect 12440 1056 12456 1120
rect 12520 1056 12528 1120
rect 12208 1055 12528 1056
<< via3 >>
rect 8216 15804 8280 15808
rect 8216 15748 8220 15804
rect 8220 15748 8276 15804
rect 8276 15748 8280 15804
rect 8216 15744 8280 15748
rect 8296 15804 8360 15808
rect 8296 15748 8300 15804
rect 8300 15748 8356 15804
rect 8356 15748 8360 15804
rect 8296 15744 8360 15748
rect 8376 15804 8440 15808
rect 8376 15748 8380 15804
rect 8380 15748 8436 15804
rect 8436 15748 8440 15804
rect 8376 15744 8440 15748
rect 8456 15804 8520 15808
rect 8456 15748 8460 15804
rect 8460 15748 8516 15804
rect 8516 15748 8520 15804
rect 8456 15744 8520 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 12216 15260 12280 15264
rect 12216 15204 12220 15260
rect 12220 15204 12276 15260
rect 12276 15204 12280 15260
rect 12216 15200 12280 15204
rect 12296 15260 12360 15264
rect 12296 15204 12300 15260
rect 12300 15204 12356 15260
rect 12356 15204 12360 15260
rect 12296 15200 12360 15204
rect 12376 15260 12440 15264
rect 12376 15204 12380 15260
rect 12380 15204 12436 15260
rect 12436 15204 12440 15260
rect 12376 15200 12440 15204
rect 12456 15260 12520 15264
rect 12456 15204 12460 15260
rect 12460 15204 12516 15260
rect 12516 15204 12520 15260
rect 12456 15200 12520 15204
rect 8216 14716 8280 14720
rect 8216 14660 8220 14716
rect 8220 14660 8276 14716
rect 8276 14660 8280 14716
rect 8216 14656 8280 14660
rect 8296 14716 8360 14720
rect 8296 14660 8300 14716
rect 8300 14660 8356 14716
rect 8356 14660 8360 14716
rect 8296 14656 8360 14660
rect 8376 14716 8440 14720
rect 8376 14660 8380 14716
rect 8380 14660 8436 14716
rect 8436 14660 8440 14716
rect 8376 14656 8440 14660
rect 8456 14716 8520 14720
rect 8456 14660 8460 14716
rect 8460 14660 8516 14716
rect 8516 14660 8520 14716
rect 8456 14656 8520 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 12216 14172 12280 14176
rect 12216 14116 12220 14172
rect 12220 14116 12276 14172
rect 12276 14116 12280 14172
rect 12216 14112 12280 14116
rect 12296 14172 12360 14176
rect 12296 14116 12300 14172
rect 12300 14116 12356 14172
rect 12356 14116 12360 14172
rect 12296 14112 12360 14116
rect 12376 14172 12440 14176
rect 12376 14116 12380 14172
rect 12380 14116 12436 14172
rect 12436 14116 12440 14172
rect 12376 14112 12440 14116
rect 12456 14172 12520 14176
rect 12456 14116 12460 14172
rect 12460 14116 12516 14172
rect 12516 14116 12520 14172
rect 12456 14112 12520 14116
rect 8216 13628 8280 13632
rect 8216 13572 8220 13628
rect 8220 13572 8276 13628
rect 8276 13572 8280 13628
rect 8216 13568 8280 13572
rect 8296 13628 8360 13632
rect 8296 13572 8300 13628
rect 8300 13572 8356 13628
rect 8356 13572 8360 13628
rect 8296 13568 8360 13572
rect 8376 13628 8440 13632
rect 8376 13572 8380 13628
rect 8380 13572 8436 13628
rect 8436 13572 8440 13628
rect 8376 13568 8440 13572
rect 8456 13628 8520 13632
rect 8456 13572 8460 13628
rect 8460 13572 8516 13628
rect 8516 13572 8520 13628
rect 8456 13568 8520 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 12216 13084 12280 13088
rect 12216 13028 12220 13084
rect 12220 13028 12276 13084
rect 12276 13028 12280 13084
rect 12216 13024 12280 13028
rect 12296 13084 12360 13088
rect 12296 13028 12300 13084
rect 12300 13028 12356 13084
rect 12356 13028 12360 13084
rect 12296 13024 12360 13028
rect 12376 13084 12440 13088
rect 12376 13028 12380 13084
rect 12380 13028 12436 13084
rect 12436 13028 12440 13084
rect 12376 13024 12440 13028
rect 12456 13084 12520 13088
rect 12456 13028 12460 13084
rect 12460 13028 12516 13084
rect 12516 13028 12520 13084
rect 12456 13024 12520 13028
rect 8216 12540 8280 12544
rect 8216 12484 8220 12540
rect 8220 12484 8276 12540
rect 8276 12484 8280 12540
rect 8216 12480 8280 12484
rect 8296 12540 8360 12544
rect 8296 12484 8300 12540
rect 8300 12484 8356 12540
rect 8356 12484 8360 12540
rect 8296 12480 8360 12484
rect 8376 12540 8440 12544
rect 8376 12484 8380 12540
rect 8380 12484 8436 12540
rect 8436 12484 8440 12540
rect 8376 12480 8440 12484
rect 8456 12540 8520 12544
rect 8456 12484 8460 12540
rect 8460 12484 8516 12540
rect 8516 12484 8520 12540
rect 8456 12480 8520 12484
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 12216 11996 12280 12000
rect 12216 11940 12220 11996
rect 12220 11940 12276 11996
rect 12276 11940 12280 11996
rect 12216 11936 12280 11940
rect 12296 11996 12360 12000
rect 12296 11940 12300 11996
rect 12300 11940 12356 11996
rect 12356 11940 12360 11996
rect 12296 11936 12360 11940
rect 12376 11996 12440 12000
rect 12376 11940 12380 11996
rect 12380 11940 12436 11996
rect 12436 11940 12440 11996
rect 12376 11936 12440 11940
rect 12456 11996 12520 12000
rect 12456 11940 12460 11996
rect 12460 11940 12516 11996
rect 12516 11940 12520 11996
rect 12456 11936 12520 11940
rect 8216 11452 8280 11456
rect 8216 11396 8220 11452
rect 8220 11396 8276 11452
rect 8276 11396 8280 11452
rect 8216 11392 8280 11396
rect 8296 11452 8360 11456
rect 8296 11396 8300 11452
rect 8300 11396 8356 11452
rect 8356 11396 8360 11452
rect 8296 11392 8360 11396
rect 8376 11452 8440 11456
rect 8376 11396 8380 11452
rect 8380 11396 8436 11452
rect 8436 11396 8440 11452
rect 8376 11392 8440 11396
rect 8456 11452 8520 11456
rect 8456 11396 8460 11452
rect 8460 11396 8516 11452
rect 8516 11396 8520 11452
rect 8456 11392 8520 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 12216 10908 12280 10912
rect 12216 10852 12220 10908
rect 12220 10852 12276 10908
rect 12276 10852 12280 10908
rect 12216 10848 12280 10852
rect 12296 10908 12360 10912
rect 12296 10852 12300 10908
rect 12300 10852 12356 10908
rect 12356 10852 12360 10908
rect 12296 10848 12360 10852
rect 12376 10908 12440 10912
rect 12376 10852 12380 10908
rect 12380 10852 12436 10908
rect 12436 10852 12440 10908
rect 12376 10848 12440 10852
rect 12456 10908 12520 10912
rect 12456 10852 12460 10908
rect 12460 10852 12516 10908
rect 12516 10852 12520 10908
rect 12456 10848 12520 10852
rect 8216 10364 8280 10368
rect 8216 10308 8220 10364
rect 8220 10308 8276 10364
rect 8276 10308 8280 10364
rect 8216 10304 8280 10308
rect 8296 10364 8360 10368
rect 8296 10308 8300 10364
rect 8300 10308 8356 10364
rect 8356 10308 8360 10364
rect 8296 10304 8360 10308
rect 8376 10364 8440 10368
rect 8376 10308 8380 10364
rect 8380 10308 8436 10364
rect 8436 10308 8440 10364
rect 8376 10304 8440 10308
rect 8456 10364 8520 10368
rect 8456 10308 8460 10364
rect 8460 10308 8516 10364
rect 8516 10308 8520 10364
rect 8456 10304 8520 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 12216 9820 12280 9824
rect 12216 9764 12220 9820
rect 12220 9764 12276 9820
rect 12276 9764 12280 9820
rect 12216 9760 12280 9764
rect 12296 9820 12360 9824
rect 12296 9764 12300 9820
rect 12300 9764 12356 9820
rect 12356 9764 12360 9820
rect 12296 9760 12360 9764
rect 12376 9820 12440 9824
rect 12376 9764 12380 9820
rect 12380 9764 12436 9820
rect 12436 9764 12440 9820
rect 12376 9760 12440 9764
rect 12456 9820 12520 9824
rect 12456 9764 12460 9820
rect 12460 9764 12516 9820
rect 12516 9764 12520 9820
rect 12456 9760 12520 9764
rect 8216 9276 8280 9280
rect 8216 9220 8220 9276
rect 8220 9220 8276 9276
rect 8276 9220 8280 9276
rect 8216 9216 8280 9220
rect 8296 9276 8360 9280
rect 8296 9220 8300 9276
rect 8300 9220 8356 9276
rect 8356 9220 8360 9276
rect 8296 9216 8360 9220
rect 8376 9276 8440 9280
rect 8376 9220 8380 9276
rect 8380 9220 8436 9276
rect 8436 9220 8440 9276
rect 8376 9216 8440 9220
rect 8456 9276 8520 9280
rect 8456 9220 8460 9276
rect 8460 9220 8516 9276
rect 8516 9220 8520 9276
rect 8456 9216 8520 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 12216 8732 12280 8736
rect 12216 8676 12220 8732
rect 12220 8676 12276 8732
rect 12276 8676 12280 8732
rect 12216 8672 12280 8676
rect 12296 8732 12360 8736
rect 12296 8676 12300 8732
rect 12300 8676 12356 8732
rect 12356 8676 12360 8732
rect 12296 8672 12360 8676
rect 12376 8732 12440 8736
rect 12376 8676 12380 8732
rect 12380 8676 12436 8732
rect 12436 8676 12440 8732
rect 12376 8672 12440 8676
rect 12456 8732 12520 8736
rect 12456 8676 12460 8732
rect 12460 8676 12516 8732
rect 12516 8676 12520 8732
rect 12456 8672 12520 8676
rect 8216 8188 8280 8192
rect 8216 8132 8220 8188
rect 8220 8132 8276 8188
rect 8276 8132 8280 8188
rect 8216 8128 8280 8132
rect 8296 8188 8360 8192
rect 8296 8132 8300 8188
rect 8300 8132 8356 8188
rect 8356 8132 8360 8188
rect 8296 8128 8360 8132
rect 8376 8188 8440 8192
rect 8376 8132 8380 8188
rect 8380 8132 8436 8188
rect 8436 8132 8440 8188
rect 8376 8128 8440 8132
rect 8456 8188 8520 8192
rect 8456 8132 8460 8188
rect 8460 8132 8516 8188
rect 8516 8132 8520 8188
rect 8456 8128 8520 8132
rect 8216 7100 8280 7104
rect 8216 7044 8220 7100
rect 8220 7044 8276 7100
rect 8276 7044 8280 7100
rect 8216 7040 8280 7044
rect 8296 7100 8360 7104
rect 8296 7044 8300 7100
rect 8300 7044 8356 7100
rect 8356 7044 8360 7100
rect 8296 7040 8360 7044
rect 8376 7100 8440 7104
rect 8376 7044 8380 7100
rect 8380 7044 8436 7100
rect 8436 7044 8440 7100
rect 8376 7040 8440 7044
rect 8456 7100 8520 7104
rect 8456 7044 8460 7100
rect 8460 7044 8516 7100
rect 8516 7044 8520 7100
rect 8456 7040 8520 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 12216 6556 12280 6560
rect 12216 6500 12220 6556
rect 12220 6500 12276 6556
rect 12276 6500 12280 6556
rect 12216 6496 12280 6500
rect 12296 6556 12360 6560
rect 12296 6500 12300 6556
rect 12300 6500 12356 6556
rect 12356 6500 12360 6556
rect 12296 6496 12360 6500
rect 12376 6556 12440 6560
rect 12376 6500 12380 6556
rect 12380 6500 12436 6556
rect 12436 6500 12440 6556
rect 12376 6496 12440 6500
rect 12456 6556 12520 6560
rect 12456 6500 12460 6556
rect 12460 6500 12516 6556
rect 12516 6500 12520 6556
rect 12456 6496 12520 6500
rect 8216 6012 8280 6016
rect 8216 5956 8220 6012
rect 8220 5956 8276 6012
rect 8276 5956 8280 6012
rect 8216 5952 8280 5956
rect 8296 6012 8360 6016
rect 8296 5956 8300 6012
rect 8300 5956 8356 6012
rect 8356 5956 8360 6012
rect 8296 5952 8360 5956
rect 8376 6012 8440 6016
rect 8376 5956 8380 6012
rect 8380 5956 8436 6012
rect 8436 5956 8440 6012
rect 8376 5952 8440 5956
rect 8456 6012 8520 6016
rect 8456 5956 8460 6012
rect 8460 5956 8516 6012
rect 8516 5956 8520 6012
rect 8456 5952 8520 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 12216 5468 12280 5472
rect 12216 5412 12220 5468
rect 12220 5412 12276 5468
rect 12276 5412 12280 5468
rect 12216 5408 12280 5412
rect 12296 5468 12360 5472
rect 12296 5412 12300 5468
rect 12300 5412 12356 5468
rect 12356 5412 12360 5468
rect 12296 5408 12360 5412
rect 12376 5468 12440 5472
rect 12376 5412 12380 5468
rect 12380 5412 12436 5468
rect 12436 5412 12440 5468
rect 12376 5408 12440 5412
rect 12456 5468 12520 5472
rect 12456 5412 12460 5468
rect 12460 5412 12516 5468
rect 12516 5412 12520 5468
rect 12456 5408 12520 5412
rect 8216 4924 8280 4928
rect 8216 4868 8220 4924
rect 8220 4868 8276 4924
rect 8276 4868 8280 4924
rect 8216 4864 8280 4868
rect 8296 4924 8360 4928
rect 8296 4868 8300 4924
rect 8300 4868 8356 4924
rect 8356 4868 8360 4924
rect 8296 4864 8360 4868
rect 8376 4924 8440 4928
rect 8376 4868 8380 4924
rect 8380 4868 8436 4924
rect 8436 4868 8440 4924
rect 8376 4864 8440 4868
rect 8456 4924 8520 4928
rect 8456 4868 8460 4924
rect 8460 4868 8516 4924
rect 8516 4868 8520 4924
rect 8456 4864 8520 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 12216 4380 12280 4384
rect 12216 4324 12220 4380
rect 12220 4324 12276 4380
rect 12276 4324 12280 4380
rect 12216 4320 12280 4324
rect 12296 4380 12360 4384
rect 12296 4324 12300 4380
rect 12300 4324 12356 4380
rect 12356 4324 12360 4380
rect 12296 4320 12360 4324
rect 12376 4380 12440 4384
rect 12376 4324 12380 4380
rect 12380 4324 12436 4380
rect 12436 4324 12440 4380
rect 12376 4320 12440 4324
rect 12456 4380 12520 4384
rect 12456 4324 12460 4380
rect 12460 4324 12516 4380
rect 12516 4324 12520 4380
rect 12456 4320 12520 4324
rect 8216 3836 8280 3840
rect 8216 3780 8220 3836
rect 8220 3780 8276 3836
rect 8276 3780 8280 3836
rect 8216 3776 8280 3780
rect 8296 3836 8360 3840
rect 8296 3780 8300 3836
rect 8300 3780 8356 3836
rect 8356 3780 8360 3836
rect 8296 3776 8360 3780
rect 8376 3836 8440 3840
rect 8376 3780 8380 3836
rect 8380 3780 8436 3836
rect 8436 3780 8440 3836
rect 8376 3776 8440 3780
rect 8456 3836 8520 3840
rect 8456 3780 8460 3836
rect 8460 3780 8516 3836
rect 8516 3780 8520 3836
rect 8456 3776 8520 3780
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 12216 3292 12280 3296
rect 12216 3236 12220 3292
rect 12220 3236 12276 3292
rect 12276 3236 12280 3292
rect 12216 3232 12280 3236
rect 12296 3292 12360 3296
rect 12296 3236 12300 3292
rect 12300 3236 12356 3292
rect 12356 3236 12360 3292
rect 12296 3232 12360 3236
rect 12376 3292 12440 3296
rect 12376 3236 12380 3292
rect 12380 3236 12436 3292
rect 12436 3236 12440 3292
rect 12376 3232 12440 3236
rect 12456 3292 12520 3296
rect 12456 3236 12460 3292
rect 12460 3236 12516 3292
rect 12516 3236 12520 3292
rect 12456 3232 12520 3236
rect 8216 2748 8280 2752
rect 8216 2692 8220 2748
rect 8220 2692 8276 2748
rect 8276 2692 8280 2748
rect 8216 2688 8280 2692
rect 8296 2748 8360 2752
rect 8296 2692 8300 2748
rect 8300 2692 8356 2748
rect 8356 2692 8360 2748
rect 8296 2688 8360 2692
rect 8376 2748 8440 2752
rect 8376 2692 8380 2748
rect 8380 2692 8436 2748
rect 8436 2692 8440 2748
rect 8376 2688 8440 2692
rect 8456 2748 8520 2752
rect 8456 2692 8460 2748
rect 8460 2692 8516 2748
rect 8516 2692 8520 2748
rect 8456 2688 8520 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 12216 2204 12280 2208
rect 12216 2148 12220 2204
rect 12220 2148 12276 2204
rect 12276 2148 12280 2204
rect 12216 2144 12280 2148
rect 12296 2204 12360 2208
rect 12296 2148 12300 2204
rect 12300 2148 12356 2204
rect 12356 2148 12360 2204
rect 12296 2144 12360 2148
rect 12376 2204 12440 2208
rect 12376 2148 12380 2204
rect 12380 2148 12436 2204
rect 12436 2148 12440 2204
rect 12376 2144 12440 2148
rect 12456 2204 12520 2208
rect 12456 2148 12460 2204
rect 12460 2148 12516 2204
rect 12516 2148 12520 2204
rect 12456 2144 12520 2148
rect 8216 1660 8280 1664
rect 8216 1604 8220 1660
rect 8220 1604 8276 1660
rect 8276 1604 8280 1660
rect 8216 1600 8280 1604
rect 8296 1660 8360 1664
rect 8296 1604 8300 1660
rect 8300 1604 8356 1660
rect 8356 1604 8360 1660
rect 8296 1600 8360 1604
rect 8376 1660 8440 1664
rect 8376 1604 8380 1660
rect 8380 1604 8436 1660
rect 8436 1604 8440 1660
rect 8376 1600 8440 1604
rect 8456 1660 8520 1664
rect 8456 1604 8460 1660
rect 8460 1604 8516 1660
rect 8516 1604 8520 1660
rect 8456 1600 8520 1604
rect 4216 1116 4280 1120
rect 4216 1060 4220 1116
rect 4220 1060 4276 1116
rect 4276 1060 4280 1116
rect 4216 1056 4280 1060
rect 4296 1116 4360 1120
rect 4296 1060 4300 1116
rect 4300 1060 4356 1116
rect 4356 1060 4360 1116
rect 4296 1056 4360 1060
rect 4376 1116 4440 1120
rect 4376 1060 4380 1116
rect 4380 1060 4436 1116
rect 4436 1060 4440 1116
rect 4376 1056 4440 1060
rect 4456 1116 4520 1120
rect 4456 1060 4460 1116
rect 4460 1060 4516 1116
rect 4516 1060 4520 1116
rect 4456 1056 4520 1060
rect 12216 1116 12280 1120
rect 12216 1060 12220 1116
rect 12220 1060 12276 1116
rect 12276 1060 12280 1116
rect 12216 1056 12280 1060
rect 12296 1116 12360 1120
rect 12296 1060 12300 1116
rect 12300 1060 12356 1116
rect 12356 1060 12360 1116
rect 12296 1056 12360 1060
rect 12376 1116 12440 1120
rect 12376 1060 12380 1116
rect 12380 1060 12436 1116
rect 12436 1060 12440 1116
rect 12376 1056 12440 1060
rect 12456 1116 12520 1120
rect 12456 1060 12460 1116
rect 12460 1060 12516 1116
rect 12516 1060 12520 1116
rect 12456 1056 12520 1060
<< metal4 >>
rect 4208 15264 4528 15824
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 6560 4528 8672
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5472 4528 6496
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 1120 4528 2144
rect 4208 1056 4216 1120
rect 4280 1056 4296 1120
rect 4360 1056 4376 1120
rect 4440 1056 4456 1120
rect 4520 1056 4528 1120
rect 4208 1040 4528 1056
rect 8208 15808 8528 15824
rect 8208 15744 8216 15808
rect 8280 15744 8296 15808
rect 8360 15744 8376 15808
rect 8440 15744 8456 15808
rect 8520 15744 8528 15808
rect 8208 14720 8528 15744
rect 8208 14656 8216 14720
rect 8280 14656 8296 14720
rect 8360 14656 8376 14720
rect 8440 14656 8456 14720
rect 8520 14656 8528 14720
rect 8208 13632 8528 14656
rect 8208 13568 8216 13632
rect 8280 13568 8296 13632
rect 8360 13568 8376 13632
rect 8440 13568 8456 13632
rect 8520 13568 8528 13632
rect 8208 12544 8528 13568
rect 8208 12480 8216 12544
rect 8280 12480 8296 12544
rect 8360 12480 8376 12544
rect 8440 12480 8456 12544
rect 8520 12480 8528 12544
rect 8208 11456 8528 12480
rect 8208 11392 8216 11456
rect 8280 11392 8296 11456
rect 8360 11392 8376 11456
rect 8440 11392 8456 11456
rect 8520 11392 8528 11456
rect 8208 10368 8528 11392
rect 8208 10304 8216 10368
rect 8280 10304 8296 10368
rect 8360 10304 8376 10368
rect 8440 10304 8456 10368
rect 8520 10304 8528 10368
rect 8208 9280 8528 10304
rect 8208 9216 8216 9280
rect 8280 9216 8296 9280
rect 8360 9216 8376 9280
rect 8440 9216 8456 9280
rect 8520 9216 8528 9280
rect 8208 8192 8528 9216
rect 8208 8128 8216 8192
rect 8280 8128 8296 8192
rect 8360 8128 8376 8192
rect 8440 8128 8456 8192
rect 8520 8128 8528 8192
rect 8208 7104 8528 8128
rect 8208 7040 8216 7104
rect 8280 7040 8296 7104
rect 8360 7040 8376 7104
rect 8440 7040 8456 7104
rect 8520 7040 8528 7104
rect 8208 6016 8528 7040
rect 8208 5952 8216 6016
rect 8280 5952 8296 6016
rect 8360 5952 8376 6016
rect 8440 5952 8456 6016
rect 8520 5952 8528 6016
rect 8208 4928 8528 5952
rect 8208 4864 8216 4928
rect 8280 4864 8296 4928
rect 8360 4864 8376 4928
rect 8440 4864 8456 4928
rect 8520 4864 8528 4928
rect 8208 3840 8528 4864
rect 8208 3776 8216 3840
rect 8280 3776 8296 3840
rect 8360 3776 8376 3840
rect 8440 3776 8456 3840
rect 8520 3776 8528 3840
rect 8208 2752 8528 3776
rect 8208 2688 8216 2752
rect 8280 2688 8296 2752
rect 8360 2688 8376 2752
rect 8440 2688 8456 2752
rect 8520 2688 8528 2752
rect 8208 1664 8528 2688
rect 8208 1600 8216 1664
rect 8280 1600 8296 1664
rect 8360 1600 8376 1664
rect 8440 1600 8456 1664
rect 8520 1600 8528 1664
rect 8208 1040 8528 1600
rect 12208 15264 12528 15824
rect 12208 15200 12216 15264
rect 12280 15200 12296 15264
rect 12360 15200 12376 15264
rect 12440 15200 12456 15264
rect 12520 15200 12528 15264
rect 12208 14176 12528 15200
rect 12208 14112 12216 14176
rect 12280 14112 12296 14176
rect 12360 14112 12376 14176
rect 12440 14112 12456 14176
rect 12520 14112 12528 14176
rect 12208 13088 12528 14112
rect 12208 13024 12216 13088
rect 12280 13024 12296 13088
rect 12360 13024 12376 13088
rect 12440 13024 12456 13088
rect 12520 13024 12528 13088
rect 12208 12000 12528 13024
rect 12208 11936 12216 12000
rect 12280 11936 12296 12000
rect 12360 11936 12376 12000
rect 12440 11936 12456 12000
rect 12520 11936 12528 12000
rect 12208 10912 12528 11936
rect 12208 10848 12216 10912
rect 12280 10848 12296 10912
rect 12360 10848 12376 10912
rect 12440 10848 12456 10912
rect 12520 10848 12528 10912
rect 12208 9824 12528 10848
rect 12208 9760 12216 9824
rect 12280 9760 12296 9824
rect 12360 9760 12376 9824
rect 12440 9760 12456 9824
rect 12520 9760 12528 9824
rect 12208 8736 12528 9760
rect 12208 8672 12216 8736
rect 12280 8672 12296 8736
rect 12360 8672 12376 8736
rect 12440 8672 12456 8736
rect 12520 8672 12528 8736
rect 12208 6560 12528 8672
rect 12208 6496 12216 6560
rect 12280 6496 12296 6560
rect 12360 6496 12376 6560
rect 12440 6496 12456 6560
rect 12520 6496 12528 6560
rect 12208 5472 12528 6496
rect 12208 5408 12216 5472
rect 12280 5408 12296 5472
rect 12360 5408 12376 5472
rect 12440 5408 12456 5472
rect 12520 5408 12528 5472
rect 12208 4384 12528 5408
rect 12208 4320 12216 4384
rect 12280 4320 12296 4384
rect 12360 4320 12376 4384
rect 12440 4320 12456 4384
rect 12520 4320 12528 4384
rect 12208 3296 12528 4320
rect 12208 3232 12216 3296
rect 12280 3232 12296 3296
rect 12360 3232 12376 3296
rect 12440 3232 12456 3296
rect 12520 3232 12528 3296
rect 12208 2208 12528 3232
rect 12208 2144 12216 2208
rect 12280 2144 12296 2208
rect 12360 2144 12376 2208
rect 12440 2144 12456 2208
rect 12520 2144 12528 2208
rect 12208 1120 12528 2144
rect 12208 1056 12216 1120
rect 12280 1056 12296 1120
rect 12360 1056 12376 1120
rect 12440 1056 12456 1120
rect 12520 1056 12528 1120
rect 12208 1040 12528 1056
use sky130_fd_sc_hd__fill_1  FILLER_1_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 1932 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 1380 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 1380 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 1104 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1620506760
transform 1 0 1104 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 2484 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20
timestamp 1620506760
transform 1 0 2944 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _319_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 2668 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _322_
timestamp 1620506760
transform 1 0 2208 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11
timestamp 1620506760
transform 1 0 2116 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _362_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform -1 0 3956 0 1 1632
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27
timestamp 1620506760
transform 1 0 3588 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33
timestamp 1620506760
transform 1 0 4140 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _359_
timestamp 1620506760
transform 1 0 4324 0 -1 1632
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  _268_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform -1 0 4140 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _269_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform -1 0 3588 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_2  _271_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform -1 0 5152 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 3772 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_31 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 3956 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_2  _277_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 5336 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_44
timestamp 1620506760
transform 1 0 5152 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1620506760
transform 1 0 6440 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1620506760
transform 1 0 6348 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _167_
timestamp 1620506760
transform -1 0 6808 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _168_
timestamp 1620506760
transform -1 0 6808 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56
timestamp 1620506760
transform 1 0 6256 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62
timestamp 1620506760
transform 1 0 6808 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_55
timestamp 1620506760
transform 1 0 6164 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_62
timestamp 1620506760
transform 1 0 6808 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_58
timestamp 1620506760
transform 1 0 6440 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _360_
timestamp 1620506760
transform -1 0 8924 0 1 1632
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _374_
timestamp 1620506760
transform 1 0 6992 0 -1 1632
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1620506760
transform 1 0 8924 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_85
timestamp 1620506760
transform 1 0 8924 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _169_
timestamp 1620506760
transform 1 0 9108 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1620506760
transform 1 0 9108 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _307_
timestamp 1620506760
transform -1 0 9476 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1620506760
transform 1 0 9476 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _375_
timestamp 1620506760
transform -1 0 11592 0 -1 1632
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_1_90
timestamp 1620506760
transform 1 0 9384 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_103
timestamp 1620506760
transform 1 0 10580 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 10948 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_2  _194_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 9752 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _185_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 11684 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1620506760
transform 1 0 11776 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1620506760
transform 1 0 11592 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114
timestamp 1620506760
transform 1 0 11592 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_112
timestamp 1620506760
transform 1 0 11408 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _306_
timestamp 1620506760
transform -1 0 12144 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1620506760
transform 1 0 12144 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_123
timestamp 1620506760
transform 1 0 12420 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _310_
timestamp 1620506760
transform 1 0 12328 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _321_
timestamp 1620506760
transform -1 0 12880 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_125
timestamp 1620506760
transform 1 0 12604 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[3\].id.delayint0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 13064 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_128
timestamp 1620506760
transform 1 0 12880 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1620506760
transform -1 0 13892 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1620506760
transform -1 0 13892 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_133
timestamp 1620506760
transform 1 0 13340 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_133
timestamp 1620506760
transform 1 0 13340 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1620506760
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7
timestamp 1620506760
transform 1 0 1748 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _320_
timestamp 1620506760
transform 1 0 1840 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_11
timestamp 1620506760
transform 1 0 2116 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_18
timestamp 1620506760
transform 1 0 2760 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1620506760
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _190_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 2300 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_2  _191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 2944 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1620506760
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1620506760
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_38
timestamp 1620506760
transform 1 0 4600 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _183_
timestamp 1620506760
transform -1 0 4600 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__and4_2  _272_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 4968 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_50
timestamp 1620506760
transform 1 0 5704 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_56
timestamp 1620506760
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_2  _275_
timestamp 1620506760
transform 1 0 6440 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _328_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform -1 0 6256 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_67
timestamp 1620506760
transform 1 0 7268 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_77
timestamp 1620506760
transform 1 0 8188 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_84
timestamp 1620506760
transform 1 0 8832 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_87
timestamp 1620506760
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1620506760
transform 1 0 9016 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _186_
timestamp 1620506760
transform -1 0 8188 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _193_
timestamp 1620506760
transform 1 0 8372 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_2_108
timestamp 1620506760
transform 1 0 11040 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_101
timestamp 1620506760
transform 1 0 10396 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_2  _207_
timestamp 1620506760
transform 1 0 10580 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2ai_2  _206_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 9292 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_2  _371_
timestamp 1620506760
transform 1 0 11316 0 -1 2720
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1620506760
transform -1 0 13892 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_132
timestamp 1620506760
transform 1 0 13248 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1620506760
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1620506760
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_10
timestamp 1620506760
transform 1 0 2024 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _377_
timestamp 1620506760
transform -1 0 4140 0 1 2720
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_2  _202_
timestamp 1620506760
transform 1 0 1564 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_3_33
timestamp 1620506760
transform 1 0 4140 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__o2bb2a_2  _213_
timestamp 1620506760
transform -1 0 5152 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_44
timestamp 1620506760
transform 1 0 5152 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_58
timestamp 1620506760
transform 1 0 6440 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1620506760
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_53
timestamp 1620506760
transform 1 0 5980 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_2  _215_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform -1 0 7360 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _273_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform -1 0 5980 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_3_68
timestamp 1620506760
transform 1 0 7360 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_75
timestamp 1620506760
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_82
timestamp 1620506760
transform 1 0 8648 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__or2_2  _214_
timestamp 1620506760
transform 1 0 7544 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _276_
timestamp 1620506760
transform 1 0 8188 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 8832 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_3_101
timestamp 1620506760
transform 1 0 10396 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_91
timestamp 1620506760
transform 1 0 9476 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_2  _195_
timestamp 1620506760
transform -1 0 10396 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__and4_2  _226_
timestamp 1620506760
transform -1 0 11408 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _309_
timestamp 1620506760
transform -1 0 12880 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_112
timestamp 1620506760
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_123
timestamp 1620506760
transform 1 0 12420 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_128
timestamp 1620506760
transform 1 0 12880 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1620506760
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _188_
timestamp 1620506760
transform -1 0 12420 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[3\].id.delaybuf1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 13064 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1620506760
transform -1 0 13892 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_133
timestamp 1620506760
transform 1 0 13340 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1620506760
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_13
timestamp 1620506760
transform 1 0 2300 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_2  _198_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 2484 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__a22oi_2  _201_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform -1 0 2300 0 -1 3808
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_4_28
timestamp 1620506760
transform 1 0 3680 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_43
timestamp 1620506760
transform 1 0 5060 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1620506760
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1620506760
transform 1 0 3312 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_39
timestamp 1620506760
transform 1 0 4692 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_2  _200_
timestamp 1620506760
transform 1 0 3864 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_51
timestamp 1620506760
transform 1 0 5796 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_59
timestamp 1620506760
transform 1 0 6532 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_2  _218_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform -1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__or3_2  _267_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform -1 0 6532 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _274_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform -1 0 5796 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_4_75
timestamp 1620506760
transform 1 0 8004 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_2  _216_
timestamp 1620506760
transform 1 0 8188 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1620506760
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_82
timestamp 1620506760
transform 1 0 8648 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o2111ai_2  _225_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_99
timestamp 1620506760
transform 1 0 10212 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_2  _210_
timestamp 1620506760
transform -1 0 11224 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_4_110
timestamp 1620506760
transform 1 0 11224 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _372_
timestamp 1620506760
transform 1 0 11500 0 -1 3808
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1620506760
transform -1 0 13892 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_134
timestamp 1620506760
transform 1 0 13432 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1620506760
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_19
timestamp 1620506760
transform 1 0 2852 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1620506760
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_15
timestamp 1620506760
transform 1 0 2484 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_2  _197_
timestamp 1620506760
transform -1 0 3772 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_2  _204_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 1748 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_29
timestamp 1620506760
transform 1 0 3772 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _361_
timestamp 1620506760
transform -1 0 5980 0 1 3808
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1620506760
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_53
timestamp 1620506760
transform 1 0 5980 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _212_
timestamp 1620506760
transform -1 0 7176 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_5_66
timestamp 1620506760
transform 1 0 7176 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_81
timestamp 1620506760
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_2  _217_
timestamp 1620506760
transform -1 0 8556 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _219_
timestamp 1620506760
transform 1 0 8740 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_5_88
timestamp 1620506760
transform 1 0 9200 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _373_
timestamp 1620506760
transform 1 0 9476 0 1 3808
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_1  _308_
timestamp 1620506760
transform -1 0 13340 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_112
timestamp 1620506760
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_123
timestamp 1620506760
transform 1 0 12420 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_128
timestamp 1620506760
transform 1 0 12880 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _209_
timestamp 1620506760
transform 1 0 12604 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1620506760
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _187_
timestamp 1620506760
transform -1 0 12420 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1620506760
transform -1 0 13892 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_133
timestamp 1620506760
transform 1 0 13340 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _196_
timestamp 1620506760
transform -1 0 2116 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _203_
timestamp 1620506760
transform -1 0 1656 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_6
timestamp 1620506760
transform 1 0 1656 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1620506760
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_8
timestamp 1620506760
transform 1 0 1840 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _305_
timestamp 1620506760
transform 1 0 1564 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1620506760
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1620506760
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _199_
timestamp 1620506760
transform -1 0 3588 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _192_
timestamp 1620506760
transform -1 0 2760 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_6_11
timestamp 1620506760
transform 1 0 2116 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_18
timestamp 1620506760
transform 1 0 2760 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _376_
timestamp 1620506760
transform -1 0 3956 0 1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1620506760
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_38
timestamp 1620506760
transform 1 0 4600 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_31
timestamp 1620506760
transform 1 0 3956 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _363_
timestamp 1620506760
transform -1 0 6072 0 1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1620506760
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _184_
timestamp 1620506760
transform -1 0 4600 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _270_
timestamp 1620506760
transform 1 0 4784 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _180_
timestamp 1620506760
transform -1 0 6624 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_47
timestamp 1620506760
transform 1 0 5428 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_51
timestamp 1620506760
transform 1 0 5796 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_54
timestamp 1620506760
transform 1 0 6072 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1620506760
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _164_
timestamp 1620506760
transform 1 0 6808 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _166_
timestamp 1620506760
transform 1 0 6440 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_60
timestamp 1620506760
transform 1 0 6624 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_65
timestamp 1620506760
transform 1 0 7084 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_61
timestamp 1620506760
transform 1 0 6716 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _364_
timestamp 1620506760
transform 1 0 6992 0 1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_6_70
timestamp 1620506760
transform 1 0 7544 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_85
timestamp 1620506760
transform 1 0 8924 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_76
timestamp 1620506760
transform 1 0 8096 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_84
timestamp 1620506760
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _165_
timestamp 1620506760
transform 1 0 7268 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _205_
timestamp 1620506760
transform -1 0 8096 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _234_
timestamp 1620506760
transform -1 0 9936 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1620506760
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _233_
timestamp 1620506760
transform 1 0 8280 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_96
timestamp 1620506760
transform 1 0 9936 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_105
timestamp 1620506760
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _365_
timestamp 1620506760
transform 1 0 9476 0 1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1620506760
transform 1 0 10948 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _211_
timestamp 1620506760
transform -1 0 10764 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_6_110
timestamp 1620506760
transform 1 0 11224 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_122
timestamp 1620506760
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_112
timestamp 1620506760
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _358_
timestamp 1620506760
transform 1 0 11500 0 -1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1620506760
transform -1 0 11960 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1620506760
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1620506760
transform 1 0 11960 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_2  _178_
timestamp 1620506760
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1620506760
transform -1 0 13892 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1620506760
transform -1 0 13892 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_134
timestamp 1620506760
transform 1 0 13432 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_132
timestamp 1620506760
transform 1 0 13248 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1620506760
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_12
timestamp 1620506760
transform 1 0 2208 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _349_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 1380 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform -1 0 3404 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_8_43
timestamp 1620506760
transform 1 0 5060 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_30
timestamp 1620506760
transform 1 0 3864 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1620506760
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_25
timestamp 1620506760
transform 1 0 3404 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_39
timestamp 1620506760
transform 1 0 4692 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen1
timestamp 1620506760
transform 1 0 4048 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_8_47
timestamp 1620506760
transform 1 0 5428 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _378_
timestamp 1620506760
transform 1 0 5612 0 -1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 1620506760
transform -1 0 5428 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _175_
timestamp 1620506760
transform 1 0 9108 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1620506760
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_70
timestamp 1620506760
transform 1 0 7544 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_82
timestamp 1620506760
transform 1 0 8648 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_2  _266_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 7912 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1620506760
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_102
timestamp 1620506760
transform 1 0 10488 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__o22ai_2  _265_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 9568 0 -1 5984
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[4\].id.delaybuf0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform -1 0 11224 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_110
timestamp 1620506760
transform 1 0 11224 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _357_
timestamp 1620506760
transform 1 0 11408 0 -1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1620506760
transform -1 0 13892 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_133
timestamp 1620506760
transform 1 0 13340 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1620506760
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_10
timestamp 1620506760
transform 1 0 2024 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen1
timestamp 1620506760
transform 1 0 1380 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[2\].id.delayenb0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform -1 0 3864 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_9_34
timestamp 1620506760
transform 1 0 4232 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _317_
timestamp 1620506760
transform 1 0 4324 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_38
timestamp 1620506760
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_30
timestamp 1620506760
transform 1 0 3864 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _348_
timestamp 1620506760
transform 1 0 4784 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_9_49
timestamp 1620506760
transform 1 0 5612 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_58
timestamp 1620506760
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_55
timestamp 1620506760
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1620506760
transform -1 0 6164 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _262_
timestamp 1620506760
transform -1 0 7176 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1620506760
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_80
timestamp 1620506760
transform 1 0 8464 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_66
timestamp 1620506760
transform 1 0 7176 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_76
timestamp 1620506760
transform 1 0 8096 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_2  _260_
timestamp 1620506760
transform -1 0 8096 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_2  _235_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 8556 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_89
timestamp 1620506760
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_100
timestamp 1620506760
transform 1 0 10304 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_2  _237_
timestamp 1620506760
transform 1 0 10488 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_2  _264_
timestamp 1620506760
transform 1 0 9476 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _316_
timestamp 1620506760
transform -1 0 12512 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _323_
timestamp 1620506760
transform -1 0 12972 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _324_
timestamp 1620506760
transform -1 0 13432 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_119
timestamp 1620506760
transform 1 0 12052 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_124
timestamp 1620506760
transform 1 0 12512 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_129
timestamp 1620506760
transform 1 0 12972 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1620506760
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_110
timestamp 1620506760
transform 1 0 11224 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[3\].id.delaybuf0
timestamp 1620506760
transform 1 0 11684 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1620506760
transform -1 0 13892 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_134
timestamp 1620506760
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 2576 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1620506760
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1620506760
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _345_
timestamp 1620506760
transform -1 0 3588 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[2\].id.delayenb1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 1564 0 -1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_1  _315_
timestamp 1620506760
transform 1 0 3864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1620506760
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_33
timestamp 1620506760
transform 1 0 4140 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1620506760
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[4\].id.delayenb0
timestamp 1620506760
transform 1 0 4324 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_10_53
timestamp 1620506760
transform 1 0 5980 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _366_
timestamp 1620506760
transform -1 0 8096 0 -1 7072
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_10_83
timestamp 1620506760
transform 1 0 8740 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_76
timestamp 1620506760
transform 1 0 8096 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1620506760
transform 1 0 9108 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1620506760
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _258_
timestamp 1620506760
transform 1 0 8280 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_10_90
timestamp 1620506760
transform 1 0 9384 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[3\].id.delayenb0
timestamp 1620506760
transform 1 0 9660 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_10_111
timestamp 1620506760
transform 1 0 11316 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _356_
timestamp 1620506760
transform -1 0 13432 0 -1 7072
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1620506760
transform -1 0 13892 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_134
timestamp 1620506760
transform 1 0 13432 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1620506760
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1620506760
transform 1 0 1380 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_7
timestamp 1620506760
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_16
timestamp 1620506760
transform 1 0 2576 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[2\].id.delaybuf1
timestamp 1620506760
transform -1 0 1748 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen0
timestamp 1620506760
transform 1 0 1932 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[2\].id.delaybuf0
timestamp 1620506760
transform -1 0 3128 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_22
timestamp 1620506760
transform 1 0 3128 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _318_
timestamp 1620506760
transform 1 0 3404 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_28
timestamp 1620506760
transform 1 0 3680 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_41
timestamp 1620506760
transform 1 0 4876 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[4\].id.delayenb1
timestamp 1620506760
transform 1 0 3864 0 1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_1  FILLER_11_56
timestamp 1620506760
transform 1 0 6256 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1620506760
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1620506760
transform 1 0 5888 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _344_
timestamp 1620506760
transform 1 0 6440 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen0
timestamp 1620506760
transform -1 0 5888 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_11_67
timestamp 1620506760
transform 1 0 7268 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_79
timestamp 1620506760
transform 1 0 8372 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_2  _238_
timestamp 1620506760
transform 1 0 8924 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_2  _263_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 7544 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_93
timestamp 1620506760
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_101
timestamp 1620506760
transform 1 0 10396 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _224_
timestamp 1620506760
transform -1 0 10396 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen0
timestamp 1620506760
transform 1 0 10764 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_11_112
timestamp 1620506760
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_126
timestamp 1620506760
transform 1 0 12696 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1620506760
transform 1 0 12880 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1620506760
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_115
timestamp 1620506760
transform 1 0 11684 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_131
timestamp 1620506760
transform 1 0 13156 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen1
timestamp 1620506760
transform 1 0 12052 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1620506760
transform -1 0 13892 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_135
timestamp 1620506760
transform 1 0 13524 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1620506760
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1620506760
transform 1 0 1380 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[1\].id.delayenb0
timestamp 1620506760
transform 1 0 1472 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__buf_1  _327_
timestamp 1620506760
transform 1 0 3312 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_22
timestamp 1620506760
transform 1 0 3128 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1620506760
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1620506760
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_34
timestamp 1620506760
transform 1 0 4232 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_2  _261_
timestamp 1620506760
transform 1 0 4600 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[1\].id.delaybuf0
timestamp 1620506760
transform -1 0 4232 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_52
timestamp 1620506760
transform 1 0 5888 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _314_
timestamp 1620506760
transform -1 0 5888 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_47
timestamp 1620506760
transform 1 0 5428 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_64
timestamp 1620506760
transform 1 0 6992 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _351_
timestamp 1620506760
transform 1 0 6164 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_12_80
timestamp 1620506760
transform 1 0 8464 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_69
timestamp 1620506760
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _174_
timestamp 1620506760
transform 1 0 7176 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1620506760
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _259_
timestamp 1620506760
transform -1 0 8464 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_2  _249_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 9108 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_12_96
timestamp 1620506760
transform 1 0 9936 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _370_
timestamp 1620506760
transform 1 0 10212 0 -1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_12_120
timestamp 1620506760
transform 1 0 12144 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[3\].id.delayenb1
timestamp 1620506760
transform 1 0 12328 0 -1 8160
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1620506760
transform -1 0 13892 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_133
timestamp 1620506760
transform 1 0 13340 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _350_
timestamp 1620506760
transform 1 0 1380 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[2\].id.delayint0
timestamp 1620506760
transform 1 0 1840 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[4\].id.delayint0
timestamp 1620506760
transform -1 0 1656 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_6
timestamp 1620506760
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1620506760
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1620506760
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen1
timestamp 1620506760
transform -1 0 3404 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[1\].id.delaybuf1
timestamp 1620506760
transform -1 0 2576 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_12
timestamp 1620506760
transform 1 0 2208 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_11
timestamp 1620506760
transform 1 0 2116 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_16
timestamp 1620506760
transform 1 0 2576 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[1\].id.delayenb1
timestamp 1620506760
transform -1 0 3404 0 1 8160
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_3  FILLER_14_35
timestamp 1620506760
transform 1 0 4324 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_25
timestamp 1620506760
transform 1 0 3404 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _367_
timestamp 1620506760
transform 1 0 3588 0 1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1620506760
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_25
timestamp 1620506760
transform 1 0 3404 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_2  _289_
timestamp 1620506760
transform 1 0 4600 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_1  ringosc.iss.reseten0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 3864 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _313_
timestamp 1620506760
transform 1 0 5888 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_55
timestamp 1620506760
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_46
timestamp 1620506760
transform 1 0 5336 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _368_
timestamp 1620506760
transform -1 0 7452 0 -1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1620506760
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_48
timestamp 1620506760
transform 1 0 5520 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_2  _286_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 6440 0 1 8160
box -38 -48 958 592
use sky130_fd_sc_hd__o32a_2  _241_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform -1 0 8648 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _240_
timestamp 1620506760
transform 1 0 7636 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_69
timestamp 1620506760
transform 1 0 7452 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_68
timestamp 1620506760
transform 1 0 7360 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _251_
timestamp 1620506760
transform -1 0 9016 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_14_82
timestamp 1620506760
transform 1 0 8648 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_79
timestamp 1620506760
transform 1 0 8372 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__o32a_2  _245_
timestamp 1620506760
transform -1 0 9936 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1620506760
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_86
timestamp 1620506760
transform 1 0 9016 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_96
timestamp 1620506760
transform 1 0 9936 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_105
timestamp 1620506760
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_96
timestamp 1620506760
transform 1 0 9936 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_107
timestamp 1620506760
transform 1 0 10948 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _246_
timestamp 1620506760
transform 1 0 10948 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _256_
timestamp 1620506760
transform 1 0 11132 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _250_
timestamp 1620506760
transform -1 0 10764 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _247_
timestamp 1620506760
transform -1 0 9936 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _254_
timestamp 1620506760
transform 1 0 10120 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _347_
timestamp 1620506760
transform 1 0 12052 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_110
timestamp 1620506760
transform 1 0 11224 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_115
timestamp 1620506760
transform 1 0 11684 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1620506760
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 1620506760
transform 1 0 11776 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_114
timestamp 1620506760
transform 1 0 11592 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_119
timestamp 1620506760
transform 1 0 12052 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1620506760
transform 1 0 12236 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_128
timestamp 1620506760
transform 1 0 12880 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_124
timestamp 1620506760
transform 1 0 12512 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _312_
timestamp 1620506760
transform -1 0 12972 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_129
timestamp 1620506760
transform 1 0 12972 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _311_
timestamp 1620506760
transform -1 0 13340 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _325_
timestamp 1620506760
transform -1 0 13432 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1620506760
transform -1 0 13892 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1620506760
transform -1 0 13892 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_133
timestamp 1620506760
transform 1 0 13340 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_134
timestamp 1620506760
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1620506760
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_12
timestamp 1620506760
transform 1 0 2208 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_21
timestamp 1620506760
transform 1 0 3036 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[1\].id.delayint0
timestamp 1620506760
transform 1 0 2760 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _330_
timestamp 1620506760
transform 1 0 1380 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_15_28
timestamp 1620506760
transform 1 0 3680 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _181_
timestamp 1620506760
transform 1 0 3220 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp01 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 3956 0 1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_15_44
timestamp 1620506760
transform 1 0 5152 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_58
timestamp 1620506760
transform 1 0 6440 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_62
timestamp 1620506760
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1620506760
transform -1 0 6808 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1620506760
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_53
timestamp 1620506760
transform 1 0 5980 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _227_
timestamp 1620506760
transform -1 0 7452 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _302_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform -1 0 5980 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_82
timestamp 1620506760
transform 1 0 8648 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_69
timestamp 1620506760
transform 1 0 7452 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _242_
timestamp 1620506760
transform -1 0 9568 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_2  _257_
timestamp 1620506760
transform 1 0 7820 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_92
timestamp 1620506760
transform 1 0 9568 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_102
timestamp 1620506760
transform 1 0 10488 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_2  _255_
timestamp 1620506760
transform -1 0 11316 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _243_
timestamp 1620506760
transform -1 0 10488 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_111
timestamp 1620506760
transform 1 0 11316 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_118
timestamp 1620506760
transform 1 0 11960 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_130
timestamp 1620506760
transform 1 0 13064 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _171_
timestamp 1620506760
transform -1 0 11960 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1620506760
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _339_
timestamp 1620506760
transform 1 0 12236 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1620506760
transform -1 0 13892 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1620506760
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_21
timestamp 1620506760
transform 1 0 3036 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[11\].id.delayenb0
timestamp 1620506760
transform 1 0 1380 0 -1 10336
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_16_39
timestamp 1620506760
transform 1 0 4692 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1620506760
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1620506760
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_35
timestamp 1620506760
transform 1 0 4324 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _182_
timestamp 1620506760
transform -1 0 4324 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_2  _287_
timestamp 1620506760
transform 1 0 4784 0 -1 10336
box -38 -48 958 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform -1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_54
timestamp 1620506760
transform 1 0 6072 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_65
timestamp 1620506760
transform 1 0 7084 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_50
timestamp 1620506760
transform 1 0 5704 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_2  _300_
timestamp 1620506760
transform 1 0 6164 0 -1 10336
box -38 -48 958 592
use sky130_fd_sc_hd__decap_3  FILLER_16_83
timestamp 1620506760
transform 1 0 8740 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_76
timestamp 1620506760
transform 1 0 8096 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1620506760
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _239_
timestamp 1620506760
transform 1 0 8280 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _252_
timestamp 1620506760
transform -1 0 9752 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_2  _298_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 7268 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_94
timestamp 1620506760
transform 1 0 9752 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_99
timestamp 1620506760
transform 1 0 10212 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _369_
timestamp 1620506760
transform 1 0 10396 0 -1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  _170_
timestamp 1620506760
transform 1 0 9936 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_122
timestamp 1620506760
transform 1 0 12328 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_131
timestamp 1620506760
transform 1 0 13156 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen1
timestamp 1620506760
transform 1 0 12512 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1620506760
transform -1 0 13892 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_135
timestamp 1620506760
transform 1 0 13524 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1620506760
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_6
timestamp 1620506760
transform 1 0 1656 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_15
timestamp 1620506760
transform 1 0 2484 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_20
timestamp 1620506760
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[11\].id.delayint0
timestamp 1620506760
transform -1 0 1656 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[11\].id.delaybuf1
timestamp 1620506760
transform -1 0 2944 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen0
timestamp 1620506760
transform 1 0 1840 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_17_40
timestamp 1620506760
transform 1 0 4784 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__einvn_8  ringosc.iss.delayenb0
timestamp 1620506760
transform 1 0 3128 0 1 10336
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  FILLER_17_54
timestamp 1620506760
transform 1 0 6072 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1620506760
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_58
timestamp 1620506760
transform 1 0 6440 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_2  _303_
timestamp 1620506760
transform -1 0 6072 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _297_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 6808 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_17_76
timestamp 1620506760
transform 1 0 8096 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_69
timestamp 1620506760
transform 1 0 7452 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__or2_2  _221_
timestamp 1620506760
transform 1 0 7636 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _223_
timestamp 1620506760
transform 1 0 8648 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_88
timestamp 1620506760
transform 1 0 9200 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_95
timestamp 1620506760
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_104
timestamp 1620506760
transform 1 0 10672 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__or2_2  _280_
timestamp 1620506760
transform 1 0 9384 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_2  _290_
timestamp 1620506760
transform -1 0 10672 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _299_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 10856 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_112
timestamp 1620506760
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1620506760
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_2  _292_
timestamp 1620506760
transform 1 0 11684 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1620506760
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[7\].id.delayenb1
timestamp 1620506760
transform 1 0 12328 0 1 10336
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1620506760
transform -1 0 13892 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_133
timestamp 1620506760
transform 1 0 13340 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1620506760
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_18
timestamp 1620506760
transform 1 0 2760 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1620506760
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen1
timestamp 1620506760
transform -1 0 3588 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[11\].id.delayenb1
timestamp 1620506760
transform 1 0 1748 0 -1 11424
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1620506760
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_37
timestamp 1620506760
transform 1 0 4508 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_42
timestamp 1620506760
transform 1 0 4968 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1620506760
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[4\].id.delaybuf1
timestamp 1620506760
transform 1 0 4692 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen1
timestamp 1620506760
transform -1 0 4508 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_18_51
timestamp 1620506760
transform 1 0 5796 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_56
timestamp 1620506760
transform 1 0 6256 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _172_
timestamp 1620506760
transform 1 0 5980 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_2  _295_
timestamp 1620506760
transform 1 0 6440 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_2  _284_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform -1 0 5796 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_18_80
timestamp 1620506760
transform 1 0 8464 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1620506760
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_67
timestamp 1620506760
transform 1 0 7268 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_87
timestamp 1620506760
transform 1 0 9108 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _355_
timestamp 1620506760
transform 1 0 7636 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_101
timestamp 1620506760
transform 1 0 10396 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _329_
timestamp 1620506760
transform 1 0 10580 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__o41a_2  _285_
timestamp 1620506760
transform 1 0 9476 0 -1 11424
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_18_112
timestamp 1620506760
transform 1 0 11408 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[7\].id.delayenb0
timestamp 1620506760
transform 1 0 11776 0 -1 11424
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1620506760
transform -1 0 13892 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_134
timestamp 1620506760
transform 1 0 13432 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1620506760
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1620506760
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3
timestamp 1620506760
transform 1 0 1380 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_16
timestamp 1620506760
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1620506760
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  ringosc.iss.ctrlen0
timestamp 1620506760
transform -1 0 3220 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _331_
timestamp 1620506760
transform 1 0 1748 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[10\].id.delayenb0
timestamp 1620506760
transform 1 0 1472 0 -1 12512
box -38 -48 1694 592
use sky130_fd_sc_hd__mux2_1  _354_
timestamp 1620506760
transform 1 0 3864 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.iss.delaybuf0
timestamp 1620506760
transform -1 0 3588 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1620506760
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_23
timestamp 1620506760
transform 1 0 3220 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_22
timestamp 1620506760
transform 1 0 3128 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1620506760
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  ringosc.iss.const1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 4600 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _282_
timestamp 1620506760
transform 1 0 4876 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _291_
timestamp 1620506760
transform 1 0 5060 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_19_36
timestamp 1620506760
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_41
timestamp 1620506760
transform 1 0 4876 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_39
timestamp 1620506760
transform 1 0 4692 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_4  ringosc.iss.delayenb1
timestamp 1620506760
transform 1 0 3404 0 1 11424
box -38 -48 1050 592
use sky130_fd_sc_hd__o31a_2  _283_
timestamp 1620506760
transform 1 0 5796 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_1  ringosc.iss.delayint0
timestamp 1620506760
transform 1 0 5888 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_50
timestamp 1620506760
transform 1 0 5704 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_49
timestamp 1620506760
transform 1 0 5612 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__o41a_2  _296_
timestamp 1620506760
transform 1 0 6440 0 1 11424
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1620506760
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _173_
timestamp 1620506760
transform 1 0 6716 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_55
timestamp 1620506760
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_59
timestamp 1620506760
transform 1 0 6532 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_64
timestamp 1620506760
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__o311a_2  _293_
timestamp 1620506760
transform 1 0 7176 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_2  _304_
timestamp 1620506760
transform 1 0 7912 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_75
timestamp 1620506760
transform 1 0 8004 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_68
timestamp 1620506760
transform 1 0 7360 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _294_
timestamp 1620506760
transform -1 0 8740 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_83
timestamp 1620506760
transform 1 0 8740 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_83
timestamp 1620506760
transform 1 0 8740 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1620506760
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_87
timestamp 1620506760
transform 1 0 9108 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_87
timestamp 1620506760
transform 1 0 9108 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__o31a_2  _281_
timestamp 1620506760
transform -1 0 9936 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _343_
timestamp 1620506760
transform 1 0 9292 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_96
timestamp 1620506760
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_2  _301_
timestamp 1620506760
transform -1 0 11224 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _231_
timestamp 1620506760
transform 1 0 10120 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _278_
timestamp 1620506760
transform 1 0 10304 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_20_105
timestamp 1620506760
transform 1 0 10764 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_103
timestamp 1620506760
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_98
timestamp 1620506760
transform 1 0 10120 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen1
timestamp 1620506760
transform 1 0 11132 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_19_124
timestamp 1620506760
transform 1 0 12512 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_116
timestamp 1620506760
transform 1 0 11776 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_127
timestamp 1620506760
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1620506760
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_110
timestamp 1620506760
transform 1 0 11224 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _336_
timestamp 1620506760
transform 1 0 11684 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _338_
timestamp 1620506760
transform 1 0 11960 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen0
timestamp 1620506760
transform 1 0 12696 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[8\].id.delaybuf0
timestamp 1620506760
transform -1 0 13340 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1620506760
transform -1 0 13892 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1620506760
transform -1 0 13892 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_133
timestamp 1620506760
transform 1 0 13340 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_133
timestamp 1620506760
transform 1 0 13340 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1620506760
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_12
timestamp 1620506760
transform 1 0 2208 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_21
timestamp 1620506760
transform 1 0 3036 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _332_
timestamp 1620506760
transform -1 0 2208 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen0
timestamp 1620506760
transform 1 0 2392 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_21_25
timestamp 1620506760
transform 1 0 3404 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_42
timestamp 1620506760
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_33
timestamp 1620506760
transform 1 0 4140 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _279_
timestamp 1620506760
transform -1 0 4968 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen0
timestamp 1620506760
transform 1 0 3496 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_21_58
timestamp 1620506760
transform 1 0 6440 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1620506760
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_53
timestamp 1620506760
transform 1 0 5980 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _337_
timestamp 1620506760
transform -1 0 7452 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _340_
timestamp 1620506760
transform -1 0 5980 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_69
timestamp 1620506760
transform 1 0 7452 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_74
timestamp 1620506760
transform 1 0 7912 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_81
timestamp 1620506760
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1620506760
transform 1 0 7636 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _232_
timestamp 1620506760
transform -1 0 8556 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _346_
timestamp 1620506760
transform -1 0 9568 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_92
timestamp 1620506760
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_103
timestamp 1620506760
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _335_
timestamp 1620506760
transform 1 0 9752 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen0
timestamp 1620506760
transform 1 0 10764 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_21_112
timestamp 1620506760
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1620506760
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[8\].id.delayenb0
timestamp 1620506760
transform 1 0 11684 0 1 12512
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1620506760
transform -1 0 13892 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_133
timestamp 1620506760
transform 1 0 13340 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1620506760
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1620506760
transform 1 0 1380 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_7
timestamp 1620506760
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_16
timestamp 1620506760
transform 1 0 2576 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[10\].id.delayint0
timestamp 1620506760
transform -1 0 1748 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen1
timestamp 1620506760
transform 1 0 1932 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[11\].id.delaybuf0
timestamp 1620506760
transform -1 0 3128 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_39
timestamp 1620506760
transform 1 0 4692 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _326_
timestamp 1620506760
transform -1 0 4140 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_22
timestamp 1620506760
transform 1 0 3128 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1620506760
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_33
timestamp 1620506760
transform 1 0 4140 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1620506760
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _288_
timestamp 1620506760
transform -1 0 5428 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[10\].id.delaybuf1
timestamp 1620506760
transform 1 0 3312 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[0\].id.delaybuf0
timestamp 1620506760
transform 1 0 4324 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_54
timestamp 1620506760
transform 1 0 6072 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_47
timestamp 1620506760
transform 1 0 5428 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__or2_2  _229_
timestamp 1620506760
transform -1 0 6072 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[5\].id.delayenb1
timestamp 1620506760
transform -1 0 7636 0 -1 13600
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_3  FILLER_22_83
timestamp 1620506760
transform 1 0 8740 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_71
timestamp 1620506760
transform 1 0 7636 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_77
timestamp 1620506760
transform 1 0 8188 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1620506760
transform 1 0 9108 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1620506760
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[5\].id.delaybuf0
timestamp 1620506760
transform -1 0 8188 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[6\].id.delaybuf0
timestamp 1620506760
transform 1 0 8372 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_107
timestamp 1620506760
transform 1 0 10948 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_90
timestamp 1620506760
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_103
timestamp 1620506760
transform 1 0 10580 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[8\].id.delayenb1
timestamp 1620506760
transform 1 0 11040 0 -1 13600
box -38 -48 1050 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[9\].id.delayenb1
timestamp 1620506760
transform 1 0 9568 0 -1 13600
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_6  FILLER_22_119
timestamp 1620506760
transform 1 0 12052 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_129
timestamp 1620506760
transform 1 0 12972 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[7\].id.delaybuf1
timestamp 1620506760
transform 1 0 13156 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[7\].id.delaybuf0
timestamp 1620506760
transform 1 0 12604 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1620506760
transform -1 0 13892 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_134
timestamp 1620506760
transform 1 0 13432 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1620506760
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1620506760
transform 1 0 1748 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1620506760
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_19
timestamp 1620506760
transform 1 0 2852 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[10\].id.delayenb1
timestamp 1620506760
transform 1 0 1840 0 1 13600
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_1  FILLER_23_23
timestamp 1620506760
transform 1 0 3220 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_42
timestamp 1620506760
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[0\].id.delayenb0
timestamp 1620506760
transform 1 0 3312 0 1 13600
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1620506760
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_53
timestamp 1620506760
transform 1 0 5980 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_65
timestamp 1620506760
transform 1 0 7084 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _342_
timestamp 1620506760
transform -1 0 5980 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen0
timestamp 1620506760
transform 1 0 6440 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_23_69
timestamp 1620506760
transform 1 0 7452 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[6\].id.delayenb0
timestamp 1620506760
transform 1 0 7544 0 1 13600
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  FILLER_23_88
timestamp 1620506760
transform 1 0 9200 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_98
timestamp 1620506760
transform 1 0 10120 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_107
timestamp 1620506760
transform 1 0 10948 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[8\].id.delayint0
timestamp 1620506760
transform -1 0 11408 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen0
timestamp 1620506760
transform 1 0 9476 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen1
timestamp 1620506760
transform 1 0 10304 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_23_128
timestamp 1620506760
transform 1 0 12880 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_112
timestamp 1620506760
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_119
timestamp 1620506760
transform 1 0 12052 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1620506760
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_124
timestamp 1620506760
transform 1 0 12512 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[7\].id.delayint0
timestamp 1620506760
transform 1 0 12972 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[8\].id.delaybuf1
timestamp 1620506760
transform 1 0 12236 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[9\].id.delaybuf0
timestamp 1620506760
transform -1 0 12052 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1620506760
transform -1 0 13892 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_132
timestamp 1620506760
transform 1 0 13248 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1620506760
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1620506760
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_16
timestamp 1620506760
transform 1 0 2576 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _333_
timestamp 1620506760
transform 1 0 1748 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[10\].id.delaybuf0
timestamp 1620506760
transform -1 0 3312 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_28
timestamp 1620506760
transform 1 0 3680 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_37
timestamp 1620506760
transform 1 0 4508 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1620506760
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1620506760
transform 1 0 3312 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen0
timestamp 1620506760
transform -1 0 4508 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen1
timestamp 1620506760
transform 1 0 4692 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_24_46
timestamp 1620506760
transform 1 0 5336 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[5\].id.delayenb0
timestamp 1620506760
transform 1 0 5520 0 -1 14688
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_24_87
timestamp 1620506760
transform 1 0 9108 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_66
timestamp 1620506760
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_75
timestamp 1620506760
transform 1 0 8004 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_84
timestamp 1620506760
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1620506760
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen1
timestamp 1620506760
transform -1 0 8004 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen0
timestamp 1620506760
transform 1 0 8188 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_24_106
timestamp 1620506760
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[6\].id.delayint0
timestamp 1620506760
transform 1 0 11040 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[9\].id.delayenb0
timestamp 1620506760
transform 1 0 9200 0 -1 14688
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_24_128
timestamp 1620506760
transform 1 0 12880 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_111
timestamp 1620506760
transform 1 0 11316 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[9\].id.delaybuf1
timestamp 1620506760
transform 1 0 11500 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_116 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620506760
transform 1 0 11776 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1620506760
transform -1 0 13892 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1620506760
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1620506760
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1620506760
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_27
timestamp 1620506760
transform 1 0 3588 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_40
timestamp 1620506760
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[0\].id.delayenb1
timestamp 1620506760
transform 1 0 3772 0 1 14688
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp11
timestamp 1620506760
transform -1 0 6164 0 1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_25_58
timestamp 1620506760
transform 1 0 6440 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_55
timestamp 1620506760
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1620506760
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _352_
timestamp 1620506760
transform 1 0 6716 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_25_70
timestamp 1620506760
transform 1 0 7544 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_84
timestamp 1620506760
transform 1 0 8832 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[6\].id.delayenb1
timestamp 1620506760
transform 1 0 7820 0 1 14688
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_25_99
timestamp 1620506760
transform 1 0 10212 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _334_
timestamp 1620506760
transform 1 0 9384 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _341_
timestamp 1620506760
transform 1 0 10580 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_25_127
timestamp 1620506760
transform 1 0 12788 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_112
timestamp 1620506760
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1620506760
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_115
timestamp 1620506760
transform 1 0 11684 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1620506760
transform -1 0 13892 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_135
timestamp 1620506760
transform 1 0 13524 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1620506760
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1620506760
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1620506760
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_30
timestamp 1620506760
transform 1 0 3864 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1620506760
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_34
timestamp 1620506760
transform 1 0 4232 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1620506760
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[0\].id.delayint0
timestamp 1620506760
transform -1 0 4232 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _353_
timestamp 1620506760
transform 1 0 4416 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_26_50
timestamp 1620506760
transform 1 0 5704 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_45
timestamp 1620506760
transform 1 0 5244 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_56
timestamp 1620506760
transform 1 0 6256 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1620506760
transform 1 0 6440 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_63
timestamp 1620506760
transform 1 0 6900 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[5\].id.delayint0
timestamp 1620506760
transform -1 0 6256 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[0\].id.delaybuf1
timestamp 1620506760
transform 1 0 5428 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp10
timestamp 1620506760
transform -1 0 6900 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_74
timestamp 1620506760
transform 1 0 7912 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_86
timestamp 1620506760
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1620506760
transform 1 0 9108 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_70
timestamp 1620506760
transform 1 0 7544 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_82
timestamp 1620506760
transform 1 0 8648 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[5\].id.delaybuf1
timestamp 1620506760
transform 1 0 7268 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen1
timestamp 1620506760
transform 1 0 8004 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_26_91
timestamp 1620506760
transform 1 0 9476 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[9\].id.delayint0
timestamp 1620506760
transform -1 0 10304 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[6\].id.delaybuf1
timestamp 1620506760
transform 1 0 9200 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_100
timestamp 1620506760
transform 1 0 10304 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_129
timestamp 1620506760
transform 1 0 12972 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1620506760
transform 1 0 11776 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_112
timestamp 1620506760
transform 1 0 11408 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1620506760
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1620506760
transform -1 0 13892 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_135
timestamp 1620506760
transform 1 0 13524 0 -1 15776
box -38 -48 130 592
<< labels >>
rlabel metal2 s 5538 0 5594 800 6 clockp[0]
port 0 nsew signal tristate
rlabel metal2 s 5998 16200 6054 17000 6 clockp[1]
port 1 nsew signal tristate
rlabel metal2 s 8298 16200 8354 17000 6 dco
port 2 nsew signal input
rlabel metal2 s 11058 16200 11114 17000 6 div[0]
port 3 nsew signal input
rlabel metal3 s 14200 3408 15000 3528 6 div[1]
port 4 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 div[2]
port 5 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 div[3]
port 6 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 div[4]
port 7 nsew signal input
rlabel metal2 s 13818 16200 13874 17000 6 enable
port 8 nsew signal input
rlabel metal2 s 6918 16200 6974 17000 6 ext_trim[0]
port 9 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 ext_trim[10]
port 10 nsew signal input
rlabel metal2 s 478 0 534 800 6 ext_trim[11]
port 11 nsew signal input
rlabel metal2 s 3238 16200 3294 17000 6 ext_trim[12]
port 12 nsew signal input
rlabel metal2 s 4618 16200 4674 17000 6 ext_trim[13]
port 13 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 ext_trim[14]
port 14 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 ext_trim[15]
port 15 nsew signal input
rlabel metal3 s 14200 8848 15000 8968 6 ext_trim[16]
port 16 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 ext_trim[17]
port 17 nsew signal input
rlabel metal3 s 14200 1368 15000 1488 6 ext_trim[18]
port 18 nsew signal input
rlabel metal2 s 12438 16200 12494 17000 6 ext_trim[19]
port 19 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 ext_trim[1]
port 20 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 ext_trim[20]
port 21 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 ext_trim[21]
port 22 nsew signal input
rlabel metal3 s 14200 12928 15000 13048 6 ext_trim[22]
port 23 nsew signal input
rlabel metal2 s 1858 16200 1914 17000 6 ext_trim[23]
port 24 nsew signal input
rlabel metal2 s 478 16200 534 17000 6 ext_trim[24]
port 25 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 ext_trim[25]
port 26 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 ext_trim[2]
port 27 nsew signal input
rlabel metal2 s 9678 16200 9734 17000 6 ext_trim[3]
port 28 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 ext_trim[4]
port 29 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 ext_trim[5]
port 30 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 ext_trim[6]
port 31 nsew signal input
rlabel metal3 s 14200 10888 15000 11008 6 ext_trim[7]
port 32 nsew signal input
rlabel metal3 s 14200 4768 15000 4888 6 ext_trim[8]
port 33 nsew signal input
rlabel metal3 s 14200 14968 15000 15088 6 ext_trim[9]
port 34 nsew signal input
rlabel metal3 s 14200 6808 15000 6928 6 osc
port 35 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 resetb
port 36 nsew signal input
rlabel metal4 s 12208 1040 12528 15824 6 VPWR
port 37 nsew power bidirectional
rlabel metal4 s 4208 1040 4528 15824 6 VPWR
port 38 nsew power bidirectional
rlabel metal4 s 8208 1040 8528 15824 6 VGND
port 39 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 17000
<< end >>
