magic
tech sky130A
timestamp 1624216132
<< mvnmos >>
rect 482 -264 586 -171
<< nmoslvt >>
rect -42 -269 62 -176
<< ndiff >>
rect -42 -176 62 -126
rect -42 -317 62 -269
rect 1035 -504 1069 -500
rect 1035 -526 1041 -504
rect 1063 -526 1069 -504
rect 1035 -531 1069 -526
rect 979 -550 1012 -546
rect 979 -572 985 -550
rect 1006 -572 1012 -550
rect 979 -576 1012 -572
<< mvndiff >>
rect 482 -171 586 -121
rect 482 -312 586 -264
<< ndiffc >>
rect 1041 -526 1063 -504
rect 985 -572 1006 -550
<< psubdiff >>
rect -44 -386 69 -373
rect -44 -435 -29 -386
rect 52 -435 69 -386
rect -44 -444 69 -435
rect 480 -381 593 -368
rect 480 -430 495 -381
rect 576 -430 593 -381
rect 480 -439 593 -430
<< psubdiffcont >>
rect -29 -435 52 -386
rect 495 -430 576 -381
<< poly >>
rect 978 -100 1016 -94
rect 978 -122 986 -100
rect 1007 -122 1016 -100
rect 978 -127 1016 -122
rect -107 -269 -42 -176
rect 62 -269 125 -176
rect 417 -264 482 -171
rect 586 -264 649 -171
rect 978 -194 1016 -188
rect 978 -216 986 -194
rect 1007 -216 1016 -194
rect 978 -221 1016 -216
rect 978 -247 1016 -242
rect 978 -269 986 -247
rect 1008 -269 1016 -247
rect 978 -274 1016 -269
rect 977 -352 1015 -346
rect 977 -374 985 -352
rect 1006 -374 1015 -352
rect 977 -379 1015 -374
rect 1035 -398 1073 -393
rect 1035 -420 1043 -398
rect 1065 -420 1073 -398
rect 1035 -425 1073 -420
rect 976 -504 1014 -498
rect 976 -526 984 -504
rect 1005 -526 1014 -504
rect 976 -531 1014 -526
rect 1034 -550 1072 -545
rect 1034 -572 1042 -550
rect 1064 -572 1072 -550
rect 1034 -577 1072 -572
<< polycont >>
rect 986 -122 1007 -100
rect 986 -216 1007 -194
rect 986 -269 1008 -247
rect 985 -374 1006 -352
rect 1043 -420 1065 -398
rect 984 -526 1005 -504
rect 1042 -572 1064 -550
<< locali >>
rect 954 -122 986 -100
rect 1007 -122 1099 -100
rect 954 -216 986 -194
rect 1007 -216 1099 -194
rect 954 -269 986 -247
rect 1008 -269 1099 -247
rect -44 -386 69 -373
rect -44 -435 -29 -386
rect 52 -435 69 -386
rect -44 -444 69 -435
rect 480 -381 593 -368
rect 953 -374 985 -352
rect 1006 -374 1098 -352
rect 480 -430 495 -381
rect 576 -430 593 -381
rect 953 -420 1043 -398
rect 1065 -420 1098 -398
rect 480 -439 593 -430
rect 952 -526 984 -504
rect 1005 -526 1041 -504
rect 1063 -526 1097 -504
rect 952 -572 985 -550
rect 1006 -572 1042 -550
rect 1064 -572 1097 -550
<< labels >>
flabel space 0 -38 0 -38 0 FreeSans 160 0 0 0 Derived_layers
flabel space 0 3 0 3 0 FreeSans 160 0 0 0 Exercise_5a
flabel space 1023 -6 1023 -6 0 FreeSans 160 0 0 0 Exercise_5c
flabel space 544 3 544 3 0 FreeSans 160 0 0 0 Exercise_5b
flabel space 555 -37 555 -37 0 FreeSans 160 0 0 0 Derived_layers
flabel space 1044 -48 1044 -48 0 FreeSans 160 0 0 0 Derived_layers
<< end >>
