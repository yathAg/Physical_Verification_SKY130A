* NGSPICE file created from example_por.ext - technology: sky130A

.subckt sky130_fd_sc_hvl__buf_8 A VGND VPWR X VNB VPB
X0 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=8.4e+11p pd=8.24e+06u as=1.45875e+12p ps=1.289e+07u w=750000u l=500000u
X1 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=1.68e+12p pd=1.424e+07u as=2.9175e+12p ps=2.189e+07u w=1.5e+06u l=500000u
X3 a_45_443# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=4.2375e+11p pd=4.13e+06u as=0p ps=0u w=750000u l=500000u
X4 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X5 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X6 VGND A a_45_443# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X7 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X8 VPWR A a_45_443# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.475e+11p ps=7.13e+06u w=1.5e+06u l=500000u
X9 VPWR A a_45_443# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X10 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X11 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X12 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X13 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X14 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X15 VGND A a_45_443# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X16 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X17 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X18 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X19 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X20 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X21 a_45_443# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ a_n683_n200# a_n189_n297# a_29_n297# a_189_n200#
+ a_n901_n200# a_247_n297# a_n407_n297# a_465_n297# a_407_n200# a_n625_n297# a_683_n297#
+ a_625_n200# a_n843_n297# w_n1101_n497# a_843_n200# a_n29_n200# a_n247_n200# a_n465_n200#
X0 a_n247_n200# a_n407_n297# a_n465_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=800000u
X1 a_843_n200# a_683_n297# a_625_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=800000u
X2 a_407_n200# a_247_n297# a_189_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=800000u
X3 a_189_n200# a_29_n297# a_n29_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=800000u
X4 a_n465_n200# a_n625_n297# a_n683_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=800000u
X5 a_625_n200# a_465_n297# a_407_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X6 a_n29_n200# a_n189_n297# a_n247_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X7 a_n683_n200# a_n843_n297# a_n901_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=800000u
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_TGFUGS a_n792_n200# a_298_n200# a_516_n200# a_734_n200#
+ a_n926_n422# a_138_n288# a_n298_n288# a_80_n200# a_356_n288# a_n516_n288# a_574_n288#
+ a_n734_n288# a_n138_n200# a_n356_n200# a_n574_n200# a_n80_n288#
X0 a_80_n200# a_n80_n288# a_n138_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=800000u
X1 a_n574_n200# a_n734_n288# a_n792_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=800000u
X2 a_734_n200# a_574_n288# a_516_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=800000u
X3 a_298_n200# a_138_n288# a_80_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=800000u
X4 a_n138_n200# a_n298_n288# a_n356_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=800000u
X5 a_n356_n200# a_n516_n288# a_n574_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X6 a_516_n200# a_356_n288# a_298_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_LQJW4T c1_n3036_n2800# m3_n3136_n2900#
X0 c1_n3036_n2800# m3_n3136_n2900# sky130_fd_pr__cap_mim_m3_1 l=2.8e+07u w=3e+07u
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_PBQTMM a_2826_2300# a_n2192_n2732# a_2826_n2732#
+ a_n1034_2300# a_n2578_2300# a_n1420_2300# a_n2964_2300# a_n648_n2732# a_n648_2300#
+ a_n5280_n2732# a_n3350_n2732# a_4370_2300# a_1282_n2732# a_124_n2732# a_n1420_n2732#
+ a_124_2300# a_n4894_n2732# a_n5410_n2862# a_n2964_n2732# a_510_2300# a_n4122_2300#
+ a_n4508_n2732# a_3598_2300# a_2054_2300# a_4370_n2732# a_3984_2300# a_2440_n2732#
+ a_2440_2300# a_3984_n2732# a_n2192_2300# a_n3736_2300# a_1668_2300# a_n262_n2732#
+ a_n262_2300# a_n1034_n2732# a_5142_2300# a_n2578_n2732# a_n1806_2300# a_n4122_n2732#
+ a_n5280_2300# a_2054_n2732# a_896_n2732# a_4756_2300# a_3598_n2732# a_3212_2300#
+ a_n3736_n2732# a_1668_n2732# a_n1806_n2732# a_5142_n2732# a_896_2300# a_510_n2732#
+ a_n3350_2300# a_n4508_2300# a_n4894_2300# a_3212_n2732# a_1282_2300# a_4756_n2732#
X0 a_n4122_n2732# a_n4122_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X1 a_n3736_n2732# a_n3736_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X2 a_5142_n2732# a_5142_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X3 a_n4894_n2732# a_n4894_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X4 a_1282_n2732# a_1282_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X5 a_4756_n2732# a_4756_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X6 a_124_n2732# a_124_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X7 a_896_n2732# a_896_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X8 a_510_n2732# a_510_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X9 a_n648_n2732# a_n648_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X10 a_n5280_n2732# a_n5280_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X11 a_n4508_n2732# a_n4508_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X12 a_n1034_n2732# a_n1034_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X13 a_n2192_n2732# a_n2192_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X14 a_2054_n2732# a_2054_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X15 a_1668_n2732# a_1668_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X16 a_2440_n2732# a_2440_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X17 a_n1420_n2732# a_n1420_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X18 a_n2578_n2732# a_n2578_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X19 a_3598_n2732# a_3598_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X20 a_n1806_n2732# a_n1806_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X21 a_3212_n2732# a_3212_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X22 a_n2964_n2732# a_n2964_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X23 a_2826_n2732# a_2826_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X24 a_4370_n2732# a_4370_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X25 a_3984_n2732# a_3984_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X26 a_n3350_n2732# a_n3350_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
X27 a_n262_n2732# a_n262_2300# a_n5410_n2862# sky130_fd_pr__res_xhigh_po_0p69 l=2.3e+07u
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_3YBPVB a_n80_n297# a_80_n200# w_n338_n497# a_n138_n200#
X0 a_80_n200# a_n80_n297# a_n138_n200# w_n338_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=800000u
.ends

.subckt sky130_fd_sc_hvl__schmittbuf_1 A VGND VPWR X VNB VPB
X0 X a_117_181# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=1.9875e+11p pd=2.03e+06u as=9.478e+11p ps=4.36e+06u w=750000u l=500000u
X1 a_217_207# a_117_181# a_64_207# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=2.289e+11p pd=2.77e+06u as=1.113e+11p ps=1.37e+06u w=420000u l=500000u
X2 VPWR A a_231_463# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=1.02225e+12p pd=5.2e+06u as=4.0875e+11p ps=4.09e+06u w=750000u l=500000u
X3 VGND A a_217_207# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X4 a_78_463# VGND VNB sky130_fd_pr__res_generic_nd__hv w=290000u l=1.355e+06u
X5 a_64_207# VPWR VPB sky130_fd_pr__res_generic_pd__hv w=290000u l=3.11e+06u
X6 X a_117_181# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=3.975e+11p pd=3.53e+06u as=0p ps=0u w=1.5e+06u l=500000u
X7 a_231_463# A a_117_181# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u w=750000u l=500000u
X8 a_231_463# a_117_181# a_78_463# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u w=750000u l=500000u
X9 a_217_207# A a_117_181# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=500000u
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_YUHPXE a_n80_n297# a_80_n200# w_n338_n497# a_n138_n200#
X0 a_80_n200# a_n80_n297# a_n138_n200# w_n338_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=800000u
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC a_80_n200# a_n272_n422# a_n138_n200# a_n80_n288#
X0 a_80_n200# a_n80_n288# a_n138_n200# a_n272_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=800000u
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_L4HW4T c2_n3079_n2800# m4_n3179_n2900#
X0 c2_n3079_n2800# m4_n3179_n2900# sky130_fd_pr__cap_mim_m3_2 l=2.8e+07u w=3e+07u
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_QE2A5N a_80_n200# a_n272_n422# a_n138_n200# a_n80_n288#
X0 a_80_n200# a_n80_n288# a_n138_n200# a_n272_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=800000u
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_YEUEBV a_n792_n200# a_138_n297# a_n298_n297#
+ a_298_n200# a_356_n297# a_n516_n297# a_574_n297# a_516_n200# a_n734_n297# a_734_n200#
+ a_n80_n297# a_80_n200# a_n138_n200# a_n356_n200# a_n574_n200# w_n992_n497#
X0 a_80_n200# a_n80_n297# a_n138_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=800000u
X1 a_n574_n200# a_n734_n297# a_n792_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=800000u
X2 a_734_n200# a_574_n297# a_516_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=800000u
X3 a_298_n200# a_138_n297# a_80_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=800000u
X4 a_n138_n200# a_n298_n297# a_n356_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=800000u
X5 a_n356_n200# a_n516_n297# a_n574_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X6 a_516_n200# a_356_n297# a_298_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_YUHPBG a_n80_n297# a_80_n200# w_n338_n497# a_n138_n200#
X0 a_80_n200# a_n80_n297# a_n138_n200# w_n338_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=800000u
.ends

.subckt sky130_fd_sc_hvl__inv_8 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=1.68e+12p pd=1.424e+07u as=2.055e+12p ps=1.774e+07u w=1.5e+06u l=500000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=1.14e+12p pd=1.054e+07u as=8.4e+11p ps=8.24e+06u w=750000u l=500000u
X3 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X4 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X6 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X7 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X8 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X9 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X12 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X13 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X14 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X15 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
.ends

.subckt example_por vdd3v3 vdd1v8 vss porb_h por_l porb_l
Xsky130_fd_sc_hvl__buf_8_1 sky130_fd_sc_hvl__inv_8_0/A vss vdd1v8 porb_l vss vdd1v8
+ sky130_fd_sc_hvl__buf_8
Xsky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ_0 m1_502_7653# m1_502_7653# m1_502_7653# m1_502_7653#
+ vdd3v3 m1_502_7653# m1_502_7653# m1_502_7653# vdd3v3 m1_502_7653# m1_502_7653# m1_502_7653#
+ m1_502_7653# vdd3v3 vdd3v3 vdd3v3 m1_502_7653# vdd3v3 sky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ
Xsky130_fd_pr__nfet_g5v0d10v5_TGFUGS_0 m1_721_6815# vss m1_721_6815# vss vss m1_721_6815#
+ m1_721_6815# m1_721_6815# m1_721_6815# m1_721_6815# m1_721_6815# m1_721_6815# vss
+ m1_721_6815# vss m1_721_6815# sky130_fd_pr__nfet_g5v0d10v5_TGFUGS
Xsky130_fd_pr__cap_mim_m3_1_LQJW4T_0 sky130_fd_sc_hvl__schmittbuf_1_0/A vss sky130_fd_pr__cap_mim_m3_1_LQJW4T
Xsky130_fd_pr__res_xhigh_po_0p69_PBQTMM_0 li_7954_5813# li_2935_565# li_8339_565#
+ li_4094_5813# li_2550_5813# li_4094_5813# li_2550_5813# li_4479_565# li_4866_5813#
+ vss li_2163_565# li_9498_5813# li_6795_565# li_5251_565# li_3707_565# li_5638_5813#
+ li_619_565# vss li_2163_565# li_5638_5813# li_1006_5813# li_619_565# li_8726_5813#
+ li_7182_5813# li_9883_565# li_9498_5813# li_7567_565# li_7954_5813# li_9111_565#
+ li_3322_5813# li_1778_5813# li_7182_5813# li_5251_565# li_4866_5813# li_4479_565#
+ vss li_2935_565# li_3322_5813# li_1391_565# vss li_7567_565# li_6023_565# vdd3v3
+ li_9111_565# li_8726_5813# li_1391_565# li_6795_565# li_3707_565# vss li_6410_5813#
+ li_6023_565# li_1778_5813# li_1006_5813# vss li_8339_565# li_6410_5813# li_9883_565#
+ sky130_fd_pr__res_xhigh_po_0p69_PBQTMM
Xsky130_fd_pr__pfet_g5v0d10v5_3YBPVB_0 m1_185_6573# m1_721_6815# vdd3v3 m1_2993_7658#
+ sky130_fd_pr__pfet_g5v0d10v5_3YBPVB
Xsky130_fd_sc_hvl__schmittbuf_1_0 sky130_fd_sc_hvl__schmittbuf_1_0/A vss vdd3v3 sky130_fd_sc_hvl__inv_8_0/A
+ vss vdd3v3 sky130_fd_sc_hvl__schmittbuf_1
Xsky130_fd_pr__pfet_g5v0d10v5_3YBPVB_1 m1_2756_6794# m1_4283_8081# vdd3v3 m1_2756_6794#
+ sky130_fd_pr__pfet_g5v0d10v5_3YBPVB
Xsky130_fd_pr__pfet_g5v0d10v5_3YBPVB_2 m1_2756_6794# sky130_fd_sc_hvl__schmittbuf_1_0/A
+ vdd3v3 m1_6249_7690# sky130_fd_pr__pfet_g5v0d10v5_3YBPVB
Xsky130_fd_pr__pfet_g5v0d10v5_3YBPVB_3 m1_185_6573# m1_502_7653# vdd3v3 m1_185_6573#
+ sky130_fd_pr__pfet_g5v0d10v5_3YBPVB
Xsky130_fd_pr__pfet_g5v0d10v5_YUHPXE_0 m1_4283_8081# m1_6249_7690# vdd3v3 vdd3v3 sky130_fd_pr__pfet_g5v0d10v5_YUHPXE
Xsky130_fd_pr__nfet_g5v0d10v5_ZK8HQC_1 m1_185_6573# vss vss li_2550_5813# sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC
Xsky130_fd_pr__cap_mim_m3_2_L4HW4T_0 vss sky130_fd_sc_hvl__schmittbuf_1_0/A sky130_fd_pr__cap_mim_m3_2_L4HW4T
Xsky130_fd_pr__nfet_g5v0d10v5_QE2A5N_0 m1_2756_6794# vss vss m1_721_6815# sky130_fd_pr__nfet_g5v0d10v5_QE2A5N
Xsky130_fd_pr__pfet_g5v0d10v5_YEUEBV_0 vdd3v3 m1_4283_8081# m1_4283_8081# m1_4283_8081#
+ m1_4283_8081# m1_4283_8081# m1_4283_8081# vdd3v3 m1_4283_8081# m1_4283_8081# m1_4283_8081#
+ vdd3v3 m1_4283_8081# vdd3v3 m1_4283_8081# vdd3v3 sky130_fd_pr__pfet_g5v0d10v5_YEUEBV
Xsky130_fd_pr__pfet_g5v0d10v5_YUHPBG_0 m1_502_7653# m1_2993_7658# vdd3v3 vdd3v3 sky130_fd_pr__pfet_g5v0d10v5_YUHPBG
Xsky130_fd_sc_hvl__inv_8_0 sky130_fd_sc_hvl__inv_8_0/A vss vdd1v8 por_l vss vdd1v8
+ sky130_fd_sc_hvl__inv_8
Xsky130_fd_sc_hvl__buf_8_0 sky130_fd_sc_hvl__inv_8_0/A vss vdd3v3 porb_h vss vdd3v3
+ sky130_fd_sc_hvl__buf_8
.ends

