magic
tech sky130A
magscale 1 2
timestamp 1665642826
<< locali >>
rect -642 -1132 -322 1876
rect -44 -178 24 -164
rect -44 -214 -28 -178
rect 10 -214 24 -178
rect -44 -228 24 -214
rect 334 -166 528 -142
rect 334 -322 362 -166
rect 502 -322 528 -166
rect 334 -344 528 -322
rect -642 -1440 -636 -1132
rect -328 -1440 -322 -1132
rect -642 -1446 -322 -1440
<< viali >>
rect -28 -214 10 -178
rect 362 -322 502 -166
rect 900 -224 968 -156
rect -636 -1440 -328 -1132
<< metal1 >>
rect -44 -178 24 -164
rect -44 -214 -28 -178
rect 10 -214 24 -178
rect -44 -228 24 -214
rect 334 -166 528 -142
rect 334 -322 362 -166
rect 502 -322 528 -166
rect 888 -156 980 -150
rect 888 -224 900 -156
rect 968 -224 980 -156
rect 888 -230 980 -224
rect 334 -344 528 -322
rect 1488 -477 1558 -166
rect 1482 -547 1488 -477
rect 1558 -547 1564 -477
rect -648 -1132 3044 -1126
rect -648 -1440 -636 -1132
rect -328 -1440 3044 -1132
rect -648 -1446 3044 -1440
rect 3364 -1446 3370 -1126
<< via1 >>
rect 1488 -547 1558 -477
rect 3044 -1446 3364 -1126
<< metal2 >>
rect 653 2020 963 2024
rect 648 2015 3364 2020
rect 648 1705 653 2015
rect 963 1705 3364 2015
rect 648 1700 3364 1705
rect 653 1696 963 1700
rect 1488 -477 1558 -471
rect 1871 -477 1941 -468
rect 1558 -547 1871 -477
rect 1488 -553 1558 -547
rect 1871 -556 1941 -547
rect 3044 -1126 3364 1700
rect 3044 -1452 3364 -1446
<< via2 >>
rect 653 1705 963 2015
rect 1871 -547 1941 -477
<< metal3 >>
rect 648 2015 968 2020
rect 648 1705 653 2015
rect 963 1705 968 2015
rect 648 973 968 1705
rect 648 655 649 973
rect 967 655 968 973
rect 648 654 968 655
rect 649 649 967 654
rect 1866 -172 1872 -104
rect 1940 -172 1946 -104
rect 1872 -472 1940 -172
rect 1866 -477 1946 -472
rect 1866 -547 1871 -477
rect 1941 -547 1946 -477
rect 1866 -552 1946 -547
<< via3 >>
rect 649 655 967 973
rect 1872 -172 1940 -104
<< metal4 >>
rect 648 973 2812 974
rect 648 655 649 973
rect 967 950 2812 973
rect 967 678 2516 950
rect 2788 678 2812 950
rect 967 655 2812 678
rect 648 654 2812 655
rect 1871 -104 1941 -103
rect 1871 -172 1872 -104
rect 1940 -172 2492 -104
rect 1871 -173 1941 -172
<< via4 >>
rect 2516 678 2788 950
rect 2492 -298 2812 22
<< metal5 >>
rect 2492 950 2812 974
rect 2492 678 2516 950
rect 2788 678 2812 950
rect 2492 46 2812 678
rect 2468 22 2836 46
rect 2468 -298 2492 22
rect 2812 -298 2836 22
rect 2468 -322 2836 -298
<< labels >>
flabel space -32 16 -32 16 0 FreeSans 320 0 0 0 Exercise_2a
flabel space -14 -74 -14 -74 0 FreeSans 320 0 0 0 Via_size
flabel space 438 -66 438 -66 0 FreeSans 320 0 0 0 Multiple_vias
flabel space 440 14 440 14 0 FreeSans 320 0 0 0 Exercise_2b
flabel space 1534 -66 1534 -66 0 FreeSans 320 0 0 0 Auto_generate_via
flabel space 1540 -4 1540 -4 0 FreeSans 320 0 0 0 Exercise_2d
flabel space 938 -68 938 -68 0 FreeSans 320 0 0 0 Via_overlap
flabel space 948 4 948 4 0 FreeSans 320 0 0 0 Exercise_2c
<< end >>
