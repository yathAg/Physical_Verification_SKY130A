magic
tech sky130A
magscale 1 2
timestamp 1665482633
<< error_s >>
rect -58 1876 284 1932
rect 188 1648 564 1700
rect -58 1548 382 1602
rect 116 1080 290 1082
rect 144 1052 318 1054
rect 116 970 137 1040
rect 144 1002 165 1052
rect 144 998 261 1002
rect 351 998 453 1002
rect 187 970 233 974
rect 379 970 425 974
<< pwell >>
rect -184 1932 -116 1934
rect -184 1876 284 1932
rect -184 1604 -116 1876
rect 188 1648 658 1700
rect -186 1602 -116 1604
rect -186 1548 382 1602
rect -186 1546 -116 1548
rect -186 1144 -128 1546
rect -186 1080 290 1144
rect -186 1072 -128 1080
rect -184 732 -130 1072
rect 604 998 656 1648
rect 192 762 572 808
rect -186 676 386 732
rect 498 594 570 762
<< metal1 >>
rect 196 2302 396 2402
rect -58 1994 566 2302
rect -184 1932 -116 1934
rect -184 1876 284 1932
rect -184 1604 -116 1876
rect 188 1648 658 1700
rect -186 1602 -116 1604
rect -186 1548 382 1602
rect -186 1546 -116 1548
rect -186 1450 -128 1546
rect 604 1462 656 1648
rect -506 1250 -128 1450
rect 598 1262 1028 1462
rect 598 1258 968 1262
rect -504 1246 -128 1250
rect -186 1144 -128 1246
rect -186 1080 290 1144
rect -186 1072 -128 1080
rect -184 732 -130 1072
rect 604 1054 656 1258
rect 144 998 656 1054
rect 192 762 572 808
rect -186 676 386 732
rect 498 638 570 762
rect -52 330 572 638
rect 134 208 334 330
use sky130_fd_pr__nfet_01v8_RV7F6E  XM1
timestamp 1665480844
transform 1 0 258 0 1 907
box -311 -360 311 360
use sky130_fd_pr__pfet_01v8_6LLYWG  XM2
timestamp 1665480844
transform 1 0 253 0 1 1743
box -311 -319 311 319
<< labels >>
flabel metal1 -506 1250 -306 1450 0 FreeSans 256 0 0 0 vin
port 0 nsew
flabel metal1 196 2202 396 2402 0 FreeSans 256 0 0 0 vdd
port 2 nsew
flabel metal1 828 1262 1028 1462 0 FreeSans 256 0 0 0 vout
port 3 nsew
flabel metal1 134 208 334 408 0 FreeSans 256 0 0 0 vss
port 1 nsew
<< end >>
