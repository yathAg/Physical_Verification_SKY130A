magic
tech sky130A
magscale 1 2
timestamp 1625449512
<< metal1 >>
rect -1882 138630 138118 140630
rect -1882 2630 118 138630
rect 136118 2630 138118 138630
rect -1882 642 138118 2630
rect 98 630 138118 642
<< metal2 >>
rect 2118 69960 62508 136630
rect 65092 69960 134118 136630
rect 2118 4630 62508 67680
rect 65092 4630 134118 67680
<< labels >>
flabel metal2 30492 121830 30492 121830 0 FreeSans 48000 0 0 0 Density_rules
flabel metal2 28691 132255 28691 132255 0 FreeSans 48000 0 0 0 Exercise_11
<< end >>
