magic
tech sky130A
magscale 1 2
timestamp 1665736700
<< metal1 >>
rect -220 -298 228 -258
rect -228 -488 220 -448
use sky130_fd_io__signal_5_sym_hv_local_5term  sky130_fd_io__signal_5_sym_hv_local_5term_0
timestamp 1665736700
transform 1 0 888 0 1 -2514
box 0 0 1591 2424
use sky130_fd_pr__esd_rf_nfet_20v0_hbm_21vW60p00  sky130_fd_pr__esd_rf_nfet_20v0_hbm_21vW60p00_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1665736700
transform 1 0 4132 0 1 -7360
box -1234 -1208 1534 7208
use sky130_fd_pr__nfet_01v8_EDB9KC  sky130_fd_pr__nfet_01v8_EDB9KC_0 Physical_Verification_SKY130A/Lab3_drc/paramcells
timestamp 1624216583
transform 1 0 3 0 1 -372
box -211 -252 211 252
<< labels >>
flabel space -20 42 -20 42 0 FreeSans 320 0 0 0 Exercise_6a
flabel space -12 -34 -12 -34 0 FreeSans 320 0 0 0 Parameterized_devices
flabel space 1628 50 1628 50 0 FreeSans 320 0 0 0 Exercise_6b
flabel space 1632 -34 1632 -34 0 FreeSans 320 0 0 0 PDK_devices
flabel space 4238 64 4238 64 0 FreeSans 320 0 0 0 Exercise_6c
flabel space 4220 -6 4220 -6 0 FreeSans 320 0 0 0 PDK_devices
<< end >>
