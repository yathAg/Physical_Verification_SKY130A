magic
tech sky130A
magscale 1 2
timestamp 1665861865
<< pwell >>
rect -308 -458 308 458
<< mvnmos >>
rect -80 -200 80 200
<< mvndiff >>
rect -138 188 -80 200
rect -138 -188 -126 188
rect -92 -188 -80 188
rect -138 -200 -80 -188
rect 80 188 138 200
rect 80 -188 92 188
rect 126 -188 138 188
rect 80 -200 138 -188
<< mvndiffc >>
rect -126 -188 -92 188
rect 92 -188 126 188
<< mvpsubdiff >>
rect -272 410 272 422
rect -272 376 -164 410
rect 164 376 272 410
rect -272 364 272 376
rect -272 -364 -214 364
rect 214 314 272 364
rect 214 -314 226 314
rect 260 -314 272 314
rect 214 -364 272 -314
rect -272 -376 272 -364
rect -272 -410 -164 -376
rect 164 -410 272 -376
rect -272 -422 272 -410
<< mvpsubdiffcont >>
rect -164 376 164 410
rect 226 -314 260 314
rect -164 -410 164 -376
<< poly >>
rect -80 272 80 288
rect -80 238 -64 272
rect 64 238 80 272
rect -80 200 80 238
rect -80 -238 80 -200
rect -80 -272 -64 -238
rect 64 -272 80 -238
rect -80 -288 80 -272
<< polycont >>
rect -64 238 64 272
rect -64 -272 64 -238
<< locali >>
rect -260 376 -164 410
rect 164 376 260 410
rect -260 -38 -226 376
rect 226 314 260 376
rect -80 238 -64 272
rect 64 238 80 272
rect -126 188 -92 204
rect -126 -204 -92 -188
rect 92 188 126 204
rect 92 -204 126 -188
rect -80 -272 -64 -238
rect 64 -272 80 -238
rect 226 -376 260 -314
rect -260 -410 -164 -376
rect 164 -410 260 -376
<< viali >>
rect -64 238 64 272
rect -260 -376 -226 -38
rect -126 -171 -92 -21
rect 92 21 126 171
rect -64 -272 64 -238
<< metal1 >>
rect -76 272 76 278
rect -76 238 -64 272
rect 64 238 76 272
rect -76 232 76 238
rect 86 171 132 183
rect 86 21 92 171
rect 126 21 132 171
rect 86 9 132 21
rect -132 -21 -86 -9
rect -266 -38 -220 -26
rect -266 -376 -260 -38
rect -226 -376 -220 -38
rect -132 -171 -126 -21
rect -92 -171 -86 -21
rect -132 -183 -86 -171
rect -76 -238 76 -232
rect -76 -272 -64 -238
rect 64 -272 76 -238
rect -76 -278 76 -272
rect -266 -388 -220 -376
<< properties >>
string FIXED_BBOX -243 -393 243 393
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2.00 l 0.80 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc -40 viadrn +40 viagate 100 viagb 0 viagr 0 viagl +45 viagt 0
<< end >>
