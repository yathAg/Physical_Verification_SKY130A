magic
tech sky130A
magscale 1 2
timestamp 1625580977
<< error_s >>
rect 4367 2973 4419 3083
rect 4537 2973 4589 3083
rect 4683 2953 4735 3083
rect 4765 2953 4819 3083
rect 4849 2953 4903 3083
rect 4933 2953 4987 3083
rect 5017 2953 5069 3083
rect 5123 2953 5175 3083
rect 5205 2953 5259 3083
rect 5289 2953 5343 3083
rect 5373 2953 5427 3083
rect 5457 2953 5509 3083
rect 5749 2953 5802 3083
rect 5832 2953 5886 3083
rect 5916 2999 6003 3083
rect 6033 2999 6087 3083
rect 5916 2953 5966 2999
rect 4302 2624 7046 2869
rect 4302 2303 7414 2624
rect 9734 2270 9770 2916
rect 11658 2393 11673 2793
rect 15649 2781 15839 2793
rect 15652 2778 15836 2781
rect 15664 2408 15824 2778
rect 15652 2405 15836 2408
rect 15649 2393 15839 2405
rect 9819 2358 9825 2364
rect 9895 2358 9901 2364
rect 9813 2352 9819 2358
rect 9901 2352 9907 2358
rect 4698 2254 4704 2266
rect 4722 2226 4728 2238
rect 4367 2089 4419 2199
rect 4537 2089 4589 2199
rect 4827 2089 4879 2173
rect 4909 2089 4919 2173
rect 16079 2167 16082 3090
rect 16479 2567 16482 3087
rect 18443 2987 18465 3021
rect 18497 2987 18519 3021
rect 18463 2173 18465 2207
rect 18497 2173 18499 2207
rect 4367 1885 4419 1995
rect 4537 1885 4589 1995
rect 4643 1885 4695 1995
rect 4905 1885 4919 1995
rect 4302 1536 7046 1781
rect 11552 1779 11680 1783
rect 12748 1757 12752 1802
rect 12782 1757 12786 1802
rect 4216 1460 4250 1490
rect 4156 1400 4190 1460
rect 4216 1370 4250 1400
rect 4302 1215 7230 1536
rect 11375 1285 11450 1293
rect 11369 1279 11375 1285
rect 11450 1279 11456 1285
rect 11369 1241 11375 1247
rect 11450 1241 11456 1247
rect 11375 1235 11381 1241
rect 11444 1235 11450 1241
rect 6841 1141 6899 1147
rect 6841 1107 6853 1141
rect 12005 1140 12020 1624
rect 12039 1140 12054 1590
rect 20206 1367 20215 2507
rect 15510 1157 15548 1194
rect 6841 1101 6899 1107
rect 20231 994 20271 2531
rect 7031 937 7071 971
<< nwell >>
rect 9170 2096 15752 2547
rect 16501 1551 19993 2053
<< pwell >>
rect 9563 1321 9619 1331
<< pmos >>
rect 15664 2393 15824 2793
<< pdiff >>
rect 11658 2393 11673 2793
<< mvpsubdiff >>
rect 16538 2139 19956 2207
<< mvnsubdiff >>
rect 16567 1953 19927 1987
<< locali >>
rect 9141 3027 9283 3040
rect 9141 2942 9157 3027
rect 9269 2942 9283 3027
rect 9141 2203 9283 2942
rect 15991 3025 16234 3038
rect 15991 2864 16036 3025
rect 16217 2864 16234 3025
rect 15991 2207 16234 2864
rect 12143 2203 16234 2207
rect 9141 2187 16234 2203
rect 9141 2057 16027 2187
rect 9135 1140 9221 1931
rect 12143 1802 16027 2057
rect 12143 1757 12752 1802
rect 12782 1774 16027 1802
rect 16210 2074 16234 2187
rect 16210 1953 19929 2074
rect 16210 1774 16234 1953
rect 12782 1757 16234 1774
rect 12039 1445 16234 1590
rect 12039 1140 12320 1445
rect 9135 1072 12320 1140
rect 9135 1070 9605 1072
rect 9135 944 9148 1070
rect 9386 944 9605 1070
rect 9135 943 9605 944
rect 12051 1005 12320 1072
rect 15216 1140 16234 1445
rect 15216 1005 19960 1140
rect 12051 943 19960 1005
rect 9135 902 19960 943
<< viali >>
rect 5841 3011 5875 3045
rect 6393 2943 6427 2977
rect 9157 2942 9269 3027
rect 4737 2875 4771 2909
rect 4921 2875 4955 2909
rect 5197 2875 5231 2909
rect 5473 2875 5507 2909
rect 6117 2875 6151 2909
rect 6485 2875 6519 2909
rect 6005 2807 6039 2841
rect 5105 2739 5139 2773
rect 5197 2399 5231 2433
rect 5013 2263 5047 2297
rect 4829 2195 4863 2229
rect 16036 2864 16217 3025
rect 18292 2606 18338 2812
rect 16704 2506 16907 2553
rect 18559 2506 18896 2553
rect 19885 2435 19919 2631
rect 5565 2127 5599 2161
rect 5289 1923 5323 1957
rect 6301 1855 6335 1889
rect 6761 1855 6795 1889
rect 5105 1787 5139 1821
rect 5565 1787 5599 1821
rect 5749 1787 5783 1821
rect 6485 1787 6519 1821
rect 6669 1787 6703 1821
rect 5933 1719 5967 1753
rect 5381 1379 5415 1413
rect 6853 1107 6887 1141
rect 16027 1774 16210 2187
rect 16970 1527 17228 1586
rect 9148 944 9386 1070
rect 9605 943 12051 1072
rect 12320 1005 15216 1445
rect 17539 1436 17606 1630
rect 17750 1472 17953 1519
rect 19370 1487 19416 1648
rect 5657 835 5691 869
rect 6117 835 6151 869
rect 5473 699 5507 733
rect 5933 699 5967 733
rect 6577 699 6611 733
rect 6761 699 6795 733
rect 6669 563 6703 597
<< metal1 >>
rect 4340 3082 6908 3178
rect 5829 3045 5887 3051
rect 5829 3011 5841 3045
rect 5875 3011 5887 3045
rect 5829 3005 5887 3011
rect 9140 3027 16233 3038
rect 5844 2974 5872 3005
rect 6381 2977 6439 2983
rect 6381 2974 6393 2977
rect 4740 2946 5872 2974
rect 6120 2946 6393 2974
rect 4740 2918 4768 2946
rect 4722 2906 4728 2918
rect 4635 2878 4728 2906
rect 4722 2866 4728 2878
rect 4780 2866 4786 2918
rect 4906 2866 4912 2918
rect 4964 2866 4970 2918
rect 5090 2866 5096 2918
rect 5148 2906 5154 2918
rect 5185 2909 5243 2915
rect 5185 2906 5197 2909
rect 5148 2878 5197 2906
rect 5148 2866 5154 2878
rect 5185 2875 5197 2878
rect 5231 2906 5243 2909
rect 5274 2906 5280 2918
rect 5231 2878 5280 2906
rect 5231 2875 5243 2878
rect 5185 2869 5243 2875
rect 5274 2866 5280 2878
rect 5332 2866 5338 2918
rect 5458 2906 5464 2918
rect 5371 2878 5464 2906
rect 5458 2866 5464 2878
rect 5516 2866 5522 2918
rect 6120 2915 6148 2946
rect 6381 2943 6393 2946
rect 6427 2974 6439 2977
rect 6427 2946 6908 2974
rect 6427 2943 6439 2946
rect 6381 2937 6439 2943
rect 9140 2942 9157 3027
rect 9269 3025 16233 3027
rect 9269 3021 16036 3025
rect 9724 3012 16036 3021
rect 9724 2953 10126 3012
rect 9269 2945 10126 2953
rect 16217 2961 16233 3025
rect 16384 3004 19941 3030
rect 9269 2942 16036 2945
rect 9140 2931 16036 2942
rect 6105 2909 6163 2915
rect 6105 2875 6117 2909
rect 6151 2875 6163 2909
rect 6105 2869 6163 2875
rect 6286 2866 6292 2918
rect 6344 2906 6350 2918
rect 6473 2909 6531 2915
rect 6473 2906 6485 2909
rect 6344 2878 6485 2906
rect 6344 2866 6350 2878
rect 6473 2875 6485 2878
rect 6519 2875 6531 2909
rect 6473 2869 6531 2875
rect 4998 2730 5004 2782
rect 5056 2770 5062 2782
rect 5093 2773 5151 2779
rect 5093 2770 5105 2773
rect 5056 2742 5105 2770
rect 5056 2730 5062 2742
rect 5093 2739 5105 2742
rect 5139 2739 5151 2773
rect 5476 2770 5504 2866
rect 5993 2841 6051 2847
rect 5993 2807 6005 2841
rect 6039 2838 6051 2841
rect 6304 2838 6332 2866
rect 9318 2862 9476 2879
rect 6039 2810 6332 2838
rect 6039 2807 6051 2810
rect 5993 2801 6051 2807
rect 6562 2798 6568 2850
rect 6620 2838 6626 2850
rect 6620 2810 6908 2838
rect 6620 2798 6626 2810
rect 9318 2790 9536 2862
rect 9809 2834 9819 2896
rect 9901 2881 9918 2896
rect 9901 2837 11598 2881
rect 11929 2837 12090 2881
rect 9901 2834 9918 2837
rect 9318 2776 9382 2790
rect 5476 2742 6908 2770
rect 5093 2733 5151 2739
rect 4340 2538 6908 2634
rect 5182 2430 5188 2442
rect 5143 2402 5188 2430
rect 5182 2390 5188 2402
rect 5240 2390 5246 2442
rect 9318 2393 9413 2776
rect 9475 2393 9536 2790
rect 9621 2540 9667 2792
rect 9727 2644 11921 2780
rect 9602 2405 11637 2540
rect 4814 2322 4820 2374
rect 4872 2362 4878 2374
rect 4872 2334 5228 2362
rect 4872 2322 4878 2334
rect 4640 2254 4646 2306
rect 4698 2294 4704 2306
rect 4906 2294 4912 2306
rect 4698 2266 4912 2294
rect 4698 2254 4704 2266
rect 4906 2254 4912 2266
rect 4964 2294 4970 2306
rect 5001 2297 5059 2303
rect 5001 2294 5013 2297
rect 4964 2266 5013 2294
rect 4964 2254 4970 2266
rect 5001 2263 5013 2266
rect 5047 2263 5059 2297
rect 5001 2257 5059 2263
rect 5200 2238 5228 2334
rect 9318 2320 9536 2393
rect 9621 2349 9667 2405
rect 9809 2349 9819 2358
rect 9318 2306 9475 2320
rect 9318 2253 9382 2306
rect 9621 2305 9819 2349
rect 9809 2296 9819 2305
rect 9901 2349 9918 2358
rect 11966 2349 12044 2837
rect 12093 2410 12400 2556
rect 9901 2308 12090 2349
rect 9901 2305 12022 2308
rect 9901 2296 9918 2305
rect 12460 2253 12533 2874
rect 12799 2834 13059 2880
rect 12586 2388 12656 2787
rect 4722 2186 4728 2238
rect 4780 2226 4786 2238
rect 4817 2229 4875 2235
rect 4817 2226 4829 2229
rect 4780 2198 4829 2226
rect 4780 2186 4786 2198
rect 4817 2195 4829 2198
rect 4863 2195 4875 2229
rect 4817 2189 4875 2195
rect 5182 2186 5188 2238
rect 5240 2226 5246 2238
rect 5240 2198 5858 2226
rect 9318 2205 12533 2253
rect 5240 2186 5246 2198
rect 5553 2161 5611 2167
rect 5553 2127 5565 2161
rect 5599 2158 5611 2161
rect 5734 2158 5740 2170
rect 5599 2130 5740 2158
rect 5599 2127 5611 2130
rect 5553 2121 5611 2127
rect 5734 2118 5740 2130
rect 5792 2118 5798 2170
rect 6654 2118 6660 2170
rect 6712 2158 6718 2170
rect 6712 2130 6908 2158
rect 6712 2118 6718 2130
rect 4340 1994 6908 2090
rect 9318 2000 9382 2205
rect 12597 2096 12656 2388
rect 5277 1957 5335 1963
rect 5277 1923 5289 1957
rect 5323 1954 5335 1957
rect 5323 1926 6908 1954
rect 5323 1923 5335 1926
rect 5277 1917 5335 1923
rect 6286 1886 6292 1898
rect 6247 1858 6292 1886
rect 6286 1846 6292 1858
rect 6344 1846 6350 1898
rect 6749 1889 6807 1895
rect 6749 1886 6761 1889
rect 6396 1858 6761 1886
rect 5093 1821 5151 1827
rect 5093 1787 5105 1821
rect 5139 1818 5151 1821
rect 5182 1818 5188 1830
rect 5139 1790 5188 1818
rect 5139 1787 5151 1790
rect 5093 1781 5151 1787
rect 5182 1778 5188 1790
rect 5240 1778 5246 1830
rect 5550 1778 5556 1830
rect 5608 1778 5614 1830
rect 5734 1818 5740 1830
rect 5695 1790 5740 1818
rect 5734 1778 5740 1790
rect 5792 1818 5798 1830
rect 6396 1818 6424 1858
rect 6749 1855 6761 1858
rect 6795 1886 6807 1889
rect 6795 1858 6908 1886
rect 9285 1873 9382 2000
rect 11482 2026 12656 2096
rect 12799 2394 12881 2834
rect 13383 2833 14847 2877
rect 15183 2833 15337 2877
rect 16010 2864 16036 2931
rect 16217 2864 16234 2961
rect 16384 2905 16418 3004
rect 19902 2905 19941 3004
rect 16384 2877 19941 2905
rect 13088 2557 13125 2793
rect 13209 2624 15171 2785
rect 13066 2397 14902 2557
rect 12799 2352 12873 2394
rect 12799 2306 13058 2352
rect 13088 2349 13125 2397
rect 15226 2349 15288 2833
rect 15349 2636 15637 2781
rect 15349 2442 15362 2636
rect 12799 2253 12873 2306
rect 13088 2305 15339 2349
rect 15712 2253 15774 2864
rect 12799 2205 15774 2253
rect 6795 1855 6807 1858
rect 6749 1849 6807 1855
rect 5792 1790 6424 1818
rect 6473 1821 6531 1827
rect 5792 1778 5798 1790
rect 6473 1787 6485 1821
rect 6519 1818 6531 1821
rect 6562 1818 6568 1830
rect 6519 1790 6568 1818
rect 6519 1787 6531 1790
rect 6473 1781 6531 1787
rect 5921 1753 5979 1759
rect 5921 1719 5933 1753
rect 5967 1750 5979 1753
rect 6488 1750 6516 1781
rect 6562 1778 6568 1790
rect 6620 1778 6626 1830
rect 6657 1821 6715 1827
rect 6657 1787 6669 1821
rect 6703 1787 6715 1821
rect 6657 1781 6715 1787
rect 5967 1722 6516 1750
rect 6672 1750 6700 1781
rect 6672 1722 6908 1750
rect 5967 1719 5979 1722
rect 5921 1713 5979 1719
rect 5550 1642 5556 1694
rect 5608 1682 5614 1694
rect 6562 1682 6568 1694
rect 5608 1654 6568 1682
rect 5608 1642 5614 1654
rect 6562 1642 6568 1654
rect 6620 1682 6626 1694
rect 6672 1682 6700 1722
rect 6620 1654 6700 1682
rect 9285 1721 9363 1873
rect 11482 1826 11552 2026
rect 12799 1917 12873 2205
rect 11365 1799 11375 1826
rect 6620 1642 6626 1654
rect 4340 1450 6908 1546
rect 5369 1413 5427 1419
rect 5369 1379 5381 1413
rect 5415 1410 5427 1413
rect 5550 1410 5556 1422
rect 5415 1382 5556 1410
rect 5415 1379 5427 1382
rect 5369 1373 5427 1379
rect 5550 1370 5556 1382
rect 5608 1370 5614 1422
rect 9285 1325 9382 1721
rect 6102 1098 6108 1150
rect 6160 1098 6166 1150
rect 6841 1141 6899 1147
rect 6841 1107 6853 1141
rect 6887 1138 6899 1141
rect 6887 1110 6908 1138
rect 6887 1107 6899 1110
rect 6841 1101 6899 1107
rect 9125 1070 9401 1078
rect 4340 906 6908 1002
rect 9125 944 9148 1070
rect 9386 944 9401 1070
rect 9125 937 9401 944
rect 9125 902 9233 937
rect 9445 902 9499 1785
rect 9881 1755 11375 1799
rect 11451 1779 11552 1826
rect 11867 1826 12873 1917
rect 11680 1779 11838 1799
rect 11451 1755 11838 1779
rect 9563 1497 9734 1724
rect 11482 1704 11552 1755
rect 9821 1567 11552 1704
rect 9563 1331 11660 1497
rect 9563 1321 9734 1331
rect 9605 1078 9734 1321
rect 11729 1285 11793 1755
rect 11867 1701 11942 1826
rect 15852 1817 15923 2796
rect 16010 2187 16234 2864
rect 18286 2812 18344 2824
rect 18286 2606 18292 2812
rect 18338 2803 18344 2812
rect 19228 2803 19238 2805
rect 18338 2753 19238 2803
rect 18338 2606 18344 2753
rect 19228 2751 19238 2753
rect 19390 2751 19400 2805
rect 18286 2594 18344 2606
rect 19879 2631 19925 2643
rect 16692 2553 17439 2559
rect 16692 2506 16704 2553
rect 16907 2506 17439 2553
rect 16692 2500 17439 2506
rect 17619 2553 18908 2559
rect 17619 2506 18559 2553
rect 18896 2506 18908 2553
rect 17619 2500 18908 2506
rect 19879 2480 19885 2631
rect 19919 2480 19925 2631
rect 19843 2426 19853 2480
rect 20005 2426 20015 2480
rect 19879 2423 19925 2426
rect 11856 1325 11942 1701
rect 15507 1788 15925 1817
rect 12267 1571 15274 1594
rect 12267 1445 13431 1571
rect 14378 1445 15274 1571
rect 9881 1241 11375 1285
rect 11685 1241 11839 1285
rect 12267 1078 12320 1445
rect 9593 1072 12320 1078
rect 9593 943 9605 1072
rect 12051 1005 12320 1072
rect 15216 1283 15274 1445
rect 15507 1375 15532 1788
rect 15903 1592 15925 1788
rect 16010 1774 16027 2187
rect 16210 2076 16234 2187
rect 16379 2295 19936 2322
rect 16379 2201 16406 2295
rect 17443 2201 17718 2295
rect 19749 2201 19936 2295
rect 16379 2169 19936 2201
rect 16210 2051 19932 2076
rect 16210 1876 16271 2051
rect 17420 1876 17702 2051
rect 19850 1876 19932 2051
rect 16210 1846 19932 1876
rect 16210 1774 16234 1846
rect 19616 1845 19932 1846
rect 16010 1746 16234 1774
rect 19364 1648 19422 1660
rect 17533 1630 17612 1642
rect 15903 1586 17240 1592
rect 15903 1527 16970 1586
rect 17228 1527 17240 1586
rect 15903 1521 17240 1527
rect 15903 1375 15925 1521
rect 17529 1436 17539 1630
rect 17606 1525 17616 1630
rect 17606 1519 17965 1525
rect 17606 1472 17750 1519
rect 17953 1472 17965 1519
rect 19364 1487 19370 1648
rect 19416 1586 19422 1648
rect 19416 1517 19607 1586
rect 19772 1517 19782 1586
rect 19416 1487 19422 1517
rect 19364 1475 19422 1487
rect 17606 1466 17965 1472
rect 17606 1436 17616 1466
rect 17533 1424 17612 1436
rect 15507 1352 15925 1375
rect 15216 1194 19927 1283
rect 15216 1157 15510 1194
rect 15548 1157 19927 1194
rect 15216 1071 19927 1157
rect 15216 1005 15274 1071
rect 12051 989 15274 1005
rect 19321 1012 19816 1022
rect 12051 943 15275 989
rect 9593 937 15275 943
rect 19321 939 19333 1012
rect 19800 939 19816 1012
rect 19321 928 19816 939
rect 19321 902 19415 928
rect 5645 869 5703 875
rect 5645 835 5657 869
rect 5691 835 5703 869
rect 6102 866 6108 878
rect 6063 838 6108 866
rect 5645 829 5703 835
rect 5660 798 5688 829
rect 6102 826 6108 838
rect 6160 826 6166 878
rect 5660 770 6908 798
rect 5182 690 5188 742
rect 5240 730 5246 742
rect 5461 733 5519 739
rect 5461 730 5473 733
rect 5240 702 5473 730
rect 5240 690 5246 702
rect 5461 699 5473 702
rect 5507 730 5519 733
rect 5918 730 5924 742
rect 5507 702 5924 730
rect 5507 699 5519 702
rect 5461 693 5519 699
rect 5918 690 5924 702
rect 5976 690 5982 742
rect 6562 730 6568 742
rect 6523 702 6568 730
rect 6562 690 6568 702
rect 6620 690 6626 742
rect 6749 733 6807 739
rect 6749 699 6761 733
rect 6795 730 6807 733
rect 6795 702 6908 730
rect 6795 699 6807 702
rect 6749 693 6807 699
rect 6657 597 6715 603
rect 6657 563 6669 597
rect 6703 594 6715 597
rect 6703 566 6908 594
rect 6703 563 6715 566
rect 6657 557 6715 563
rect 4340 362 6908 458
<< via1 >>
rect 4728 2909 4780 2918
rect 4728 2875 4737 2909
rect 4737 2875 4771 2909
rect 4771 2875 4780 2909
rect 4728 2866 4780 2875
rect 4912 2909 4964 2918
rect 4912 2875 4921 2909
rect 4921 2875 4955 2909
rect 4955 2875 4964 2909
rect 4912 2866 4964 2875
rect 5096 2866 5148 2918
rect 5280 2866 5332 2918
rect 5464 2909 5516 2918
rect 5464 2875 5473 2909
rect 5473 2875 5507 2909
rect 5507 2875 5516 2909
rect 5464 2866 5516 2875
rect 9160 2953 9269 3021
rect 9269 2953 9724 3021
rect 10126 2945 16036 3012
rect 16036 2945 16193 3012
rect 6292 2866 6344 2918
rect 5004 2730 5056 2782
rect 6568 2798 6620 2850
rect 9819 2834 9901 2896
rect 5188 2433 5240 2442
rect 5188 2399 5197 2433
rect 5197 2399 5231 2433
rect 5231 2399 5240 2433
rect 5188 2390 5240 2399
rect 4820 2322 4872 2374
rect 4646 2254 4698 2306
rect 4912 2254 4964 2306
rect 9819 2296 9901 2358
rect 4728 2186 4780 2238
rect 5188 2186 5240 2238
rect 5740 2118 5792 2170
rect 6660 2118 6712 2170
rect 6292 1889 6344 1898
rect 6292 1855 6301 1889
rect 6301 1855 6335 1889
rect 6335 1855 6344 1889
rect 6292 1846 6344 1855
rect 5188 1778 5240 1830
rect 5556 1821 5608 1830
rect 5556 1787 5565 1821
rect 5565 1787 5599 1821
rect 5599 1787 5608 1821
rect 5556 1778 5608 1787
rect 5740 1821 5792 1830
rect 5740 1787 5749 1821
rect 5749 1787 5783 1821
rect 5783 1787 5792 1821
rect 16418 2905 19902 3004
rect 5740 1778 5792 1787
rect 6568 1778 6620 1830
rect 5556 1642 5608 1694
rect 6568 1642 6620 1694
rect 5556 1370 5608 1422
rect 6108 1098 6160 1150
rect 11375 1755 11451 1826
rect 19238 2751 19390 2805
rect 17439 2500 17619 2559
rect 19853 2435 19885 2480
rect 19885 2435 19919 2480
rect 19919 2435 20005 2480
rect 19853 2426 20005 2435
rect 13431 1445 14378 1571
rect 11375 1241 11450 1285
rect 13431 1022 14378 1445
rect 15532 1375 15903 1788
rect 16406 2201 17443 2295
rect 17718 2201 19749 2295
rect 16271 1876 17420 2051
rect 17702 1876 19850 2051
rect 17539 1436 17606 1630
rect 19607 1517 19772 1586
rect 19333 939 19800 1012
rect 6108 869 6160 878
rect 6108 835 6117 869
rect 6117 835 6151 869
rect 6151 835 6160 869
rect 6108 826 6160 835
rect 5188 690 5240 742
rect 5924 733 5976 742
rect 5924 699 5933 733
rect 5933 699 5967 733
rect 5967 699 5976 733
rect 5924 690 5976 699
rect 6568 733 6620 742
rect 6568 699 6577 733
rect 6577 699 6611 733
rect 6611 699 6620 733
rect 6568 690 6620 699
<< metal2 >>
rect 4728 2918 4780 2924
rect 4728 2860 4780 2866
rect 4646 2306 4698 2312
rect 4646 2248 4698 2254
rect 4658 2176 4686 2248
rect 4740 2244 4768 2860
rect 4832 2380 4860 3190
rect 4912 2918 4964 2924
rect 4912 2860 4964 2866
rect 4820 2374 4872 2380
rect 4820 2316 4872 2322
rect 4924 2312 4952 2860
rect 5016 2788 5044 3190
rect 5096 2918 5148 2924
rect 5096 2860 5148 2866
rect 5004 2782 5056 2788
rect 5004 2724 5056 2730
rect 4912 2306 4964 2312
rect 4912 2248 4964 2254
rect 4728 2238 4780 2244
rect 4728 2180 4780 2186
rect 4648 2145 4686 2176
rect 4648 282 4676 2145
rect 5108 1467 5136 2860
rect 5200 2448 5228 3190
rect 5292 2924 5320 3190
rect 5476 2924 5504 3190
rect 5280 2918 5332 2924
rect 5280 2860 5332 2866
rect 5464 2918 5516 2924
rect 5464 2860 5516 2866
rect 5188 2442 5240 2448
rect 5188 2384 5240 2390
rect 5188 2238 5240 2244
rect 5188 2180 5240 2186
rect 5200 1836 5228 2180
rect 5740 2170 5792 2176
rect 5740 2112 5792 2118
rect 5752 1836 5780 2112
rect 5188 1830 5240 1836
rect 5188 1772 5240 1778
rect 5556 1830 5608 1836
rect 5556 1772 5608 1778
rect 5740 1830 5792 1836
rect 5740 1772 5792 1778
rect 5094 1458 5150 1467
rect 5094 1393 5150 1402
rect 5200 748 5228 1772
rect 5568 1700 5596 1772
rect 5556 1694 5608 1700
rect 5556 1636 5608 1642
rect 5568 1428 5596 1636
rect 5556 1422 5608 1428
rect 5556 1364 5608 1370
rect 5922 778 5978 787
rect 5188 742 5240 748
rect 5922 713 5924 722
rect 5188 684 5240 690
rect 5976 713 5978 722
rect 5924 684 5976 690
rect 6028 282 6056 3190
rect 6292 2918 6344 2924
rect 6292 2860 6344 2866
rect 6304 1904 6332 2860
rect 6580 2856 6608 3190
rect 10085 3038 16232 3039
rect 9138 3021 16232 3038
rect 9138 2953 9160 3021
rect 9724 3013 16232 3021
rect 9138 2856 9177 2953
rect 9734 2939 9986 3013
rect 16191 3012 16232 3013
rect 16193 2945 16232 3012
rect 9734 2856 9754 2939
rect 6568 2850 6620 2856
rect 9138 2813 9754 2856
rect 9819 2896 9901 2906
rect 9819 2824 9901 2834
rect 9966 2856 9986 2939
rect 16191 2856 16232 2945
rect 16384 3004 19941 3030
rect 16384 2905 16418 3004
rect 19902 2905 19941 3004
rect 16384 2877 19941 2905
rect 6568 2792 6620 2798
rect 9829 2358 9885 2824
rect 9966 2812 16232 2856
rect 19238 2808 19390 2818
rect 19238 2738 19390 2748
rect 17439 2559 17619 2569
rect 17439 2490 17619 2500
rect 9819 2286 9901 2296
rect 16379 2295 17474 2322
rect 16379 2201 16406 2295
rect 17443 2201 17474 2295
rect 6660 2170 6712 2176
rect 16379 2169 17474 2201
rect 6660 2112 6712 2118
rect 6292 1898 6344 1904
rect 6292 1840 6344 1846
rect 6568 1830 6620 1836
rect 6672 1818 6700 2112
rect 16241 2051 17455 2076
rect 16241 1876 16271 2051
rect 17420 1876 17455 2051
rect 16241 1846 17455 1876
rect 6620 1790 6700 1818
rect 11375 1826 11451 1836
rect 6568 1772 6620 1778
rect 11375 1745 11451 1755
rect 15507 1788 15925 1817
rect 6568 1694 6620 1700
rect 6568 1636 6620 1642
rect 6108 1150 6160 1156
rect 6108 1092 6160 1098
rect 6120 884 6148 1092
rect 6108 878 6160 884
rect 6108 820 6160 826
rect 6580 748 6608 1636
rect 11388 1285 11440 1745
rect 13408 1601 14398 1620
rect 13408 1022 13431 1601
rect 14378 1022 14398 1601
rect 15507 1375 15532 1788
rect 15903 1375 15925 1788
rect 17543 1640 17600 2490
rect 19853 2483 20005 2493
rect 19853 2413 20005 2423
rect 17688 2295 19767 2322
rect 17687 2201 17718 2295
rect 19749 2201 19767 2295
rect 17688 2169 19767 2201
rect 17667 2051 19898 2076
rect 17667 1876 17702 2051
rect 19850 1876 19898 2051
rect 17667 1846 19898 1876
rect 17539 1630 17606 1640
rect 17539 1426 17606 1436
rect 15507 1352 15925 1375
rect 13408 1001 14398 1022
rect 19321 1022 19531 1846
rect 19598 1517 19607 1586
rect 19772 1517 19857 1586
rect 20009 1517 20018 1586
rect 19321 1012 19816 1022
rect 19321 939 19333 1012
rect 19800 939 19816 1012
rect 19321 928 19816 939
rect 6568 742 6620 748
rect 6568 684 6620 690
rect 4634 212 4690 282
rect 6014 212 6070 282
<< via2 >>
rect 5094 1402 5150 1458
rect 5922 742 5978 778
rect 5922 722 5924 742
rect 5924 722 5976 742
rect 5976 722 5978 742
rect 9177 2953 9724 3013
rect 9724 2953 9734 3013
rect 9177 2856 9734 2953
rect 9986 3012 16191 3013
rect 9986 2945 10126 3012
rect 10126 2945 16191 3012
rect 9986 2856 16191 2945
rect 16418 2905 19902 3004
rect 19238 2805 19390 2808
rect 19238 2751 19390 2805
rect 19238 2748 19390 2751
rect 16406 2201 17443 2295
rect 13431 1571 14378 1601
rect 13431 1274 14378 1571
rect 15532 1375 15903 1788
rect 19853 2480 20005 2483
rect 19853 2426 20005 2480
rect 19853 2423 20005 2426
rect 17718 2201 19749 2295
rect 19857 1517 20009 1586
<< metal3 >>
rect 9138 3013 16226 3035
rect 9138 2996 9177 3013
rect 9734 2996 9986 3013
rect 9138 2752 9173 2996
rect 16191 2856 16226 3013
rect 16384 3004 19941 3030
rect 16384 2905 16418 3004
rect 19902 2905 19941 3004
rect 16384 2877 19941 2905
rect 16173 2752 16226 2856
rect 9138 2717 16226 2752
rect 19228 2808 19395 2816
rect 19228 2748 19238 2808
rect 19390 2748 19531 2808
rect 19228 2743 19395 2748
rect 19471 2668 19531 2748
rect 19471 2608 20403 2668
rect 19843 2483 20010 2491
rect 19843 2423 19853 2483
rect 20005 2423 20010 2483
rect 19843 2418 20010 2423
rect 16379 2295 19767 2322
rect 16379 2201 16406 2295
rect 19749 2201 19767 2295
rect 19892 2303 19952 2418
rect 19892 2243 20404 2303
rect 16379 2169 19767 2201
rect 13211 2029 14399 2069
rect 13211 1601 13450 2029
rect 14368 1601 14399 2029
rect 4190 1460 4216 1490
rect 5089 1460 5155 1463
rect 4190 1458 5155 1460
rect 4190 1402 5094 1458
rect 5150 1402 5155 1458
rect 4190 1400 5155 1402
rect 4190 1370 4216 1400
rect 5089 1397 5155 1400
rect 13211 1274 13431 1601
rect 14378 1274 14399 1601
rect 15508 1788 15925 1817
rect 15508 1375 15532 1788
rect 15903 1375 15925 1788
rect 19847 1586 20018 1592
rect 19847 1517 19857 1586
rect 20009 1517 20402 1586
rect 19847 1510 20018 1517
rect 15508 1352 15925 1375
rect 13211 1246 14399 1274
rect 13211 1003 13407 1246
rect 5917 780 5983 783
rect 5917 778 6908 780
rect 5917 722 5922 778
rect 5978 722 6908 778
rect 5917 720 6908 722
rect 5917 717 5983 720
<< via3 >>
rect 9173 2856 9177 2996
rect 9177 2856 9734 2996
rect 9734 2856 9986 2996
rect 9986 2856 16173 2996
rect 16418 2905 19902 3004
rect 9173 2752 16173 2856
rect 16406 2201 17443 2295
rect 17443 2201 17718 2295
rect 17718 2201 19749 2295
rect 13450 1601 14368 2029
rect 13450 1310 14368 1601
rect 15532 1375 15903 1788
<< metal4 >>
rect 9138 2996 16226 3035
rect 9138 2752 9173 2996
rect 16173 2752 16226 2996
rect 9138 2717 16226 2752
rect 16341 3004 20240 3043
rect 16341 2905 16418 3004
rect 19902 2905 20240 3004
rect 16341 2714 20240 2905
rect 19943 2507 20238 2526
rect 9138 2295 19767 2407
rect 9138 2201 16406 2295
rect 19749 2201 19767 2295
rect 9138 2029 19767 2201
rect 9138 2007 13450 2029
rect 12917 1310 13450 2007
rect 14368 2007 19767 2029
rect 14368 1310 14399 2007
rect 19943 1826 19979 2507
rect 15486 1788 19979 1826
rect 15486 1375 15532 1788
rect 15903 1375 19979 1788
rect 15486 1367 19979 1375
rect 20206 1367 20238 2507
rect 15486 1343 20238 1367
rect 12917 1274 14399 1310
rect 12917 902 13111 1274
rect 13201 902 13893 1003
<< via4 >>
rect 13450 1310 14368 1999
rect 19979 1367 20206 2507
<< metal5 >>
rect 19951 2507 20231 2531
rect 13413 1999 14399 2069
rect 13413 1310 13450 1999
rect 14368 1310 14399 1999
rect 13413 1246 14399 1310
rect 13607 902 14399 1246
rect 19951 1367 19979 2507
rect 20206 1367 20231 2507
rect 19951 994 20231 1367
use sky130_fd_sc_hd__fill_1  FILLER_1_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625580977
transform 1 0 5168 0 1 954
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625580977
transform 1 0 4616 0 1 954
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625580977
transform 1 0 4340 0 1 954
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11
timestamp 1625580977
transform 1 0 5352 0 -1 954
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1625580977
transform 1 0 4340 0 -1 954
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625580977
transform 1 0 4616 0 -1 954
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625580977
transform 1 0 5720 0 -1 954
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _319_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625580977
transform 1 0 5904 0 -1 954
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20
timestamp 1625580977
transform 1 0 6180 0 -1 954
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_2  _269_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625580977
transform -1 0 6824 0 -1 954
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _322_
timestamp 1625580977
transform 1 0 5444 0 -1 954
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _362_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625580977
transform -1 0 7192 0 1 954
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625580977
transform 1 0 7002 0 -1 954
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27
timestamp 1625580977
transform 1 0 6824 0 -1 954
box -38 -48 222 592
use sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC  sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC_1 paramcells
timestamp 1625580977
transform -1 0 9471 0 1 1521
box -308 -458 308 458
use sky130_fd_pr__nfet_g5v0d10v5_TGFUGS  sky130_fd_pr__nfet_g5v0d10v5_TGFUGS_0 paramcells
timestamp 1625580977
transform 1 0 10615 0 1 1521
box -962 -458 962 458
use sky130_fd_pr__nfet_g5v0d10v5_PKVMTM  sky130_fd_pr__nfet_g5v0d10v5_PKVMTM_0 paramcells
timestamp 1625580977
transform 1 0 11760 0 1 1522
box -308 -458 308 458
use sky130_fd_sc_hvl__schmittbuf_1  sky130_fd_sc_hvl__schmittbuf_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1625580977
transform 1 0 16567 0 1 1156
box -66 -43 1122 897
use sky130_fd_sc_hvl__fill_4  sky130_fd_sc_hvl__fill_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1625580977
transform 1 0 19543 0 1 1156
box -66 -43 450 897
use sky130_fd_sc_hvl__buf_8  sky130_fd_sc_hvl__buf_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1625580977
transform 1 0 17623 0 1 1156
box -66 -43 1986 897
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1625580977
transform 1 0 4616 0 1 2042
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1625580977
transform 1 0 4340 0 1 2042
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _202_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625580977
transform 1 0 4800 0 1 2042
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_3_10
timestamp 1625580977
transform 1 0 5260 0 1 2042
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_11
timestamp 1625580977
transform 1 0 5352 0 -1 2042
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _320_
timestamp 1625580977
transform 1 0 5076 0 -1 2042
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7
timestamp 1625580977
transform 1 0 4984 0 -1 2042
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625580977
transform 1 0 4616 0 -1 2042
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1625580977
transform 1 0 4340 0 -1 2042
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_18
timestamp 1625580977
transform 1 0 5996 0 -1 2042
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_2  _191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625580977
transform 1 0 6180 0 -1 2042
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _190_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625580977
transform 1 0 5536 0 -1 2042
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_2  _377_
timestamp 1625580977
transform -1 0 7376 0 1 2042
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1625580977
transform 1 0 6824 0 -1 2042
box -38 -48 222 592
use sky130_fd_pr__pfet_g5v0d10v5_3YBPVB  sky130_fd_pr__pfet_g5v0d10v5_3YBPVB_3 paramcells
timestamp 1625580977
transform 1 0 9510 0 1 2593
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ  sky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ_0 paramcells
timestamp 1625580977
transform 1 0 10757 0 1 2593
box -1101 -497 1101 497
use sky130_fd_pr__pfet_g5v0d10v5_YUHPBG  sky130_fd_pr__pfet_g5v0d10v5_YUHPBG_0 paramcells
timestamp 1625580977
transform 1 0 12006 0 1 2593
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_3YBPVB  sky130_fd_pr__pfet_g5v0d10v5_3YBPVB_1
timestamp 1625580977
transform 1 0 12978 0 1 2593
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_3YBPVB  sky130_fd_pr__pfet_g5v0d10v5_3YBPVB_0
timestamp 1625580977
transform 1 0 12492 0 1 2593
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_YEUEBV  sky130_fd_pr__pfet_g5v0d10v5_YEUEBV_0 paramcells
timestamp 1625580977
transform 1 0 14118 0 1 2593
box -992 -497 992 497
use sky130_fd_pr__pfet_g5v0d10v5_YUHPXE  sky130_fd_pr__pfet_g5v0d10v5_YUHPXE_0 paramcells
timestamp 1625580977
transform 1 0 15258 0 1 2593
box -338 -497 338 497
use sky130_fd_sc_hvl__buf_8  sky130_fd_sc_hvl__buf_8_1
timestamp 1625580977
transform 1 0 16545 0 1 2190
box -66 -43 1986 897
use sky130_fd_pr__pfet_g5v0d10v5_3YBPVB  sky130_fd_pr__pfet_g5v0d10v5_3YBPVB_2
timestamp 1625580977
transform 1 0 15744 0 1 2593
box -338 -497 338 497
use sky130_fd_sc_hvl__inv_8  sky130_fd_sc_hvl__inv_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1625580977
transform 1 0 18497 0 1 2190
box -66 -43 1506 897
use sky130_fd_sc_hd__fill_2  FILLER_4_13
timestamp 1625580977
transform 1 0 5536 0 -1 3130
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1625580977
transform 1 0 4340 0 -1 3130
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_2  _201_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625580977
transform -1 0 5536 0 -1 3130
box -38 -48 958 592
use sky130_fd_sc_hd__a2bb2o_2  _198_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625580977
transform 1 0 5720 0 -1 3130
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1625580977
transform 1 0 6548 0 -1 3130
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_28
timestamp 1625580977
transform 1 0 6916 0 -1 3130
box -38 -48 130 592
<< labels >>
flabel metal4 s 9138 2717 9173 3035 0 FreeSans 320 0 0 0 vdd3v3
port 0 nsew
flabel metal4 s 9138 2007 9332 2407 0 FreeSans 320 0 0 0 vss
port 2 nsew
flabel metal4 s 20034 2714 20240 3043 0 FreeSans 320 0 0 0 vdd1v8
port 1 nsew
flabel metal3 20249 2243 20404 2303 0 FreeSans 320 0 0 0 por_l
port 4 nsew
flabel metal3 20248 2608 20403 2668 0 FreeSans 320 0 0 0 porb_l
port 5 nsew
flabel metal3 20029 1517 20402 1586 0 FreeSans 320 0 0 0 porb_h
port 3 nsew
<< end >>
