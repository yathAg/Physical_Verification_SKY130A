* NGSPICE file created from digital_pll.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VPWR Q VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X2 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=1.2307e+12p pd=1.144e+07u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X3 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X4 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=1.4795e+12p pd=1.507e+07u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X14 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X15 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X19 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X20 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X22 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X26 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X29 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or3_2 A B C VGND VPWR X VNB VPB
X0 VPWR a_30_53# X VPB sky130_fd_pr__pfet_01v8_hvt ad=6.115e+11p pd=5.31e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 VGND a_30_53# X VNB sky130_fd_pr__nfet_01v8 ad=5.024e+11p pd=5.23e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 X a_30_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_112_297# C a_30_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4 X a_30_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X6 a_30_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND C a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_184_297# B a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9 VPWR A a_184_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=590000u
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=1.05e+06u
.ends

.subckt sky130_fd_sc_hd__clkinv_1 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.268e+11p pd=2.22e+06u as=4.536e+11p ps=4.44e+06u w=840000u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=1.197e+11p pd=1.41e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VPWR X VNB VPB
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=4.553e+11p pd=4.29e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=5.155e+11p pd=4.31e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VPWR X VNB VPB
X0 a_79_21# C1 a_635_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=4.2e+11p ps=2.84e+06u w=1e+06u l=150000u
X1 VPWR A2 a_319_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.11e+12p pd=8.22e+06u as=7.6e+11p ps=5.52e+06u w=1e+06u l=150000u
X2 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=7.605e+11p pd=6.24e+06u as=4.355e+11p ps=3.94e+06u w=650000u l=150000u
X3 a_417_47# A2 a_319_47# VNB sky130_fd_pr__nfet_01v8 ad=2.405e+11p pd=2.04e+06u as=2.21e+11p ps=1.98e+06u w=650000u l=150000u
X4 a_79_21# A1 a_417_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_319_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X7 a_319_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X9 a_319_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_635_297# B1 a_319_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VPWR X VNB VPB
X0 VPWR a_82_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=8.098e+11p pd=7.22e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 a_646_47# B2 a_82_21# VNB sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2 a_574_369# a_313_47# a_82_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.616e+11p pd=3.69e+06u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X3 a_574_369# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 VGND a_82_21# X VNB sky130_fd_pr__nfet_01v8 ad=8.0515e+11p pd=7.55e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X5 VPWR B2 a_574_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 X a_82_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_82_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_313_47# A2_N a_313_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.696e+11p pd=1.81e+06u as=1.344e+11p ps=1.7e+06u w=640000u l=150000u
X9 a_313_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X10 a_313_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 VGND A2_N a_313_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_82_21# a_313_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND B1 a_646_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__einvp_2 A TE VGND VPWR Z VNB VPB
X0 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=4.202e+11p pd=4.22e+06u as=8.249e+11p ps=7.57e+06u w=940000u l=150000u
X1 a_204_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=5.135e+11p pd=5.48e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 VPWR TE a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X3 Z A a_204_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X5 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_204_47# TE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.63e+11p ps=3.77e+06u w=650000u l=150000u
X7 VGND TE a_204_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X9 VGND TE a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__einvn_8 A TE_B VGND VPWR Z VNB VPB
X0 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=2.3452e+12p pd=2.234e+07u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X1 VGND a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=8.71e+11p pd=9.18e+06u as=1.61525e+12p ps=1.667e+07u w=650000u l=150000u
X2 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u
X3 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.3263e+12p ps=1.231e+07u w=940000u l=150000u
X7 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X10 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X12 a_215_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_215_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_215_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X17 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X19 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X23 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X24 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X30 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_215_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 VPWR TE_B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X33 VGND TE_B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VPWR X VNB VPB
X0 X a_91_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=1.245e+12p ps=8.49e+06u w=1e+06u l=150000u
X1 a_91_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=5.35e+11p pd=5.07e+06u as=0p ps=0u w=1e+06u l=150000u
X2 a_360_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=4.6475e+11p pd=4.03e+06u as=8.8725e+11p ps=6.63e+06u w=650000u l=150000u
X3 VPWR B1 a_91_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_360_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=3.5e+11p pd=2.7e+06u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A2 a_360_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_360_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_91_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_91_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X9 X a_91_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_677_47# B1 a_360_47# VNB sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X11 a_460_297# A2 a_360_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=4.2e+11p pd=2.84e+06u as=0p ps=0u w=1e+06u l=150000u
X12 a_91_21# C1 a_677_47# VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X13 a_91_21# A3 a_460_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2_2 A B VGND VPWR X VNB VPB
X0 a_121_297# B a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1 X a_39_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=4.917e+11p ps=5.19e+06u w=650000u l=150000u
X2 VPWR a_39_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=5.715e+11p pd=5.23e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3 X a_39_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND a_39_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND A a_39_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X7 a_39_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VPWR X VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=5.63e+11p pd=5.18e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=3.6625e+11p ps=3.78e+06u w=650000u l=150000u
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__einvn_4 A TE_B VGND VPWR Z VNB VPB
X0 VGND a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=5.2e+11p pd=5.5e+06u as=9.1325e+11p ps=9.31e+06u w=650000u l=150000u
X1 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=1.2976e+12p pd=1.242e+07u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X2 VGND a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.187e+11p pd=7.47e+06u as=0p ps=0u w=940000u l=150000u
X4 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X5 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X6 a_215_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X10 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X11 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_215_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR TE_B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND TE_B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_2 A B VGND VPWR Y VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=7.9e+11p pd=7.58e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=5.135e+11p pd=5.48e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VPWR X VNB VPB
X0 VPWR a_38_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=9.2e+11p pd=7.84e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 VPWR A1 a_497_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X2 X a_38_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_141_47# B2 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X4 a_497_297# A2 a_38_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.1e+12p ps=6.2e+06u w=1e+06u l=150000u
X5 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=5.135e+11p pd=5.48e+06u as=0p ps=0u w=650000u l=150000u
X6 VPWR C1 a_38_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_237_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.25e+11p pd=2.45e+06u as=0p ps=0u w=1e+06u l=150000u
X8 a_38_47# B2 a_237_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_38_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X11 a_141_47# C1 a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.3725e+11p ps=2.03e+06u w=650000u l=150000u
X12 VGND a_38_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_225_47# B1 a_141_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_1 A VGND VPWR X VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.291e+11p pd=2.16e+06u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=1.508e+11p ps=1.62e+06u w=520000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=1.97e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=1.97e+06u
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VPWR X VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.85e+11p pd=5.17e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=2.457e+11p pd=2.85e+06u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VPWR X VNB VPB
X0 VPWR A2 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.6e+11p pd=7.72e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1 a_277_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_79_21# B1 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=0p ps=0u w=1e+06u l=150000u
X3 a_277_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=5.135e+11p pd=5.48e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X6 a_361_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X7 a_277_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.535e+11p ps=2.08e+06u w=650000u l=150000u
X9 a_79_21# A1 a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VPWR X VNB VPB
X0 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=8.45e+11p pd=7.69e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 VGND A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=5.4925e+11p pd=5.59e+06u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X2 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=1.495e+11p ps=1.76e+06u w=650000u l=150000u
X5 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.2e+11p pd=5.04e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X6 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_381_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VPWR X VNB VPB
X0 VPWR A3 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=9.6e+11p pd=7.92e+06u as=8e+11p ps=7.6e+06u w=1e+06u l=150000u
X1 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_352_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=2.3075e+11p pd=2.01e+06u as=7.5725e+11p ps=6.23e+06u w=650000u l=150000u
X3 a_549_47# A1 a_21_199# VNB sky130_fd_pr__nfet_01v8 ad=2.795e+11p pd=2.16e+06u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X4 X a_21_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=5.2e+11p pd=5.04e+06u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_21_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X6 a_665_47# A2 a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X7 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_299_297# B1 a_21_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X9 a_21_199# B2 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND A3 a_665_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR a_21_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_21_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_21_199# B1 a_352_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VPWR X VNB VPB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=2.291e+11p pd=2.16e+06u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=1.508e+11p ps=1.62e+06u w=520000u l=150000u
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VPWR Y VNB VPB
X0 VGND A2 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=4.355e+11p pd=3.94e+06u as=7.085e+11p ps=7.38e+06u w=650000u l=150000u
X1 Y B1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=8.5e+11p pd=7.7e+06u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u
X3 VPWR A1 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.3e+11p ps=5.26e+06u w=1e+06u l=150000u
X4 a_29_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A2 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND A1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_112_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_112_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_29_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_29_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_2 A B VGND VPWR Y VNB VPB
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VPWR X VNB VPB
X0 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=5.453e+11p pd=4.43e+06u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X1 VGND D a_304_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=1.1245e+12p ps=8.77e+06u w=1e+06u l=150000u
X3 a_198_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=1.596e+11p pd=1.6e+06u as=1.239e+11p ps=1.43e+06u w=420000u l=150000u
X4 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.667e+11p pd=2.95e+06u as=0p ps=0u w=420000u l=150000u
X5 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_304_47# C a_198_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VPWR X VNB VPB
X0 a_301_47# B2 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=5.85e+11p pd=5.7e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X1 VGND A2 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=5.135e+11p pd=5.48e+06u as=0p ps=0u w=650000u l=150000u
X2 a_383_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=1.34e+12p ps=8.68e+06u w=1e+06u l=150000u
X3 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X4 a_301_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X6 X a_81_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_81_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A1 a_579_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X9 a_81_21# B1 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_579_297# A2 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.7e+11p ps=2.94e+06u w=1e+06u l=150000u
X11 a_81_21# B2 a_383_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=5.2e+11p ps=5.04e+06u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VPWR X VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=8.6e+11p pd=7.72e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=5.07e+11p ps=5.46e+06u w=650000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.3e+11p pd=5.06e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X4 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=6.045e+11p ps=5.76e+06u w=650000u l=150000u
X6 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X7 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=4.73e+06u
.ends

.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VPWR Y VNB VPB
X0 VGND A2 a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=6.5975e+11p pd=5.93e+06u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.575e+11p ps=3.7e+06u w=650000u l=150000u
X2 Y A1 a_114_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X3 a_114_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=1.19e+12p pd=1.038e+07u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.5e+11p ps=5.1e+06u w=1e+06u l=150000u
X6 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_285_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=2.89e+06u
.ends

.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VPWR X VNB VPB
X0 a_108_21# B1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=3.9e+11p ps=3.8e+06u w=650000u l=150000u
X1 a_346_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.3125e+11p ps=6.15e+06u w=650000u l=150000u
X2 X a_108_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=2.275e+11p pd=2e+06u as=0p ps=0u w=650000u l=150000u
X3 a_108_21# A3 a_430_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=4.25e+11p pd=2.85e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X4 a_430_297# A2 a_346_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X5 VPWR a_108_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=1.135e+12p pd=8.27e+06u as=3.5e+11p ps=2.7e+06u w=1e+06u l=150000u
X6 a_346_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A2 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_108_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR B1 a_108_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND a_108_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_346_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VPWR Y VNB VPB
X0 Y A2 a_734_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X1 a_300_47# B2 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=9.165e+11p pd=9.32e+06u as=6.89e+11p ps=7.32e+06u w=650000u l=150000u
X2 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.685e+12p ps=1.137e+07u w=1e+06u l=150000u
X3 a_300_47# B1 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X5 a_300_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_734_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_28_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X8 Y C1 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR B1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X11 a_382_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_28_47# B1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_28_47# B2 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y B2 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR A1 a_734_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND A2 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_382_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_734_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__einvp_1 A TE VGND VPWR Z VNB VPB
X0 a_276_297# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=3.65e+11p pd=2.73e+06u as=6.415e+11p ps=3.37e+06u w=1e+06u l=150000u
X1 Z A a_204_47# VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=4.7125e+11p ps=2.75e+06u w=650000u l=150000u
X2 VPWR TE a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3 Z A a_276_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X4 a_204_47# TE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.94e+11p ps=1.95e+06u w=650000u l=150000u
X5 VGND TE a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and3_2 A B C VGND VPWR X VNB VPB
X0 VPWR a_29_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=6.749e+11p pd=6.59e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 X a_29_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.5795e+11p ps=2.99e+06u w=420000u l=150000u
X3 VGND a_29_311# X VNB sky130_fd_pr__nfet_01v8 ad=4.3955e+11p pd=4.06e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X4 a_184_53# B a_112_53# VNB sky130_fd_pr__nfet_01v8 ad=1.071e+11p pd=1.35e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X5 VPWR C a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_29_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_112_53# A a_29_311# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8 a_29_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND C a_184_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VPWR X VNB VPB
X0 VPWR A1 a_485_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.93e+11p pd=8.08e+06u as=5.3e+11p ps=5.06e+06u w=1e+06u l=150000u
X1 a_485_297# a_297_93# a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2 a_297_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=7.2375e+11p ps=7.48e+06u w=420000u l=150000u
X3 a_581_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X5 a_79_21# a_297_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A2 a_581_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X8 a_297_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_485_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VPWR X VNB VPB
X0 VGND A2 a_393_47# VNB sky130_fd_pr__nfet_01v8 ad=7.9625e+11p pd=7.65e+06u as=7.3125e+11p ps=6.15e+06u w=650000u l=150000u
X1 a_496_297# A4 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=6.05e+11p ps=3.21e+06u w=1e+06u l=150000u
X2 a_393_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A1 a_697_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.28e+12p pd=8.56e+06u as=3.5e+11p ps=2.7e+06u w=1e+06u l=150000u
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X6 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A4 a_393_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_697_297# A2 a_597_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.5e+11p ps=2.7e+06u w=1e+06u l=150000u
X9 a_393_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_393_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X12 a_597_297# A3 a_496_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VPWR X VNB VPB
X0 a_294_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=1.323e+11p pd=1.47e+06u as=4.959e+11p ps=5.21e+06u w=420000u l=150000u
X1 VPWR A2_N a_295_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.2138e+12p pd=9.74e+06u as=3.46e+11p ps=2.8e+06u w=640000u l=150000u
X2 VPWR B1 a_665_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.728e+11p ps=1.82e+06u w=640000u l=150000u
X3 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X4 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_581_47# a_295_369# a_84_21# VNB sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X7 a_665_369# B2 a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.856e+11p ps=1.86e+06u w=640000u l=150000u
X8 VGND B2 a_581_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_295_369# A2_N a_294_47# VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_84_21# a_295_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_295_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 a_581_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPB VPWR VNB
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06u area=4.347e+11p
.ends

.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VPWR X VNB VPB
X0 VPWR A1 a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.325e+12p pd=8.65e+06u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X1 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=5.4925e+11p pd=5.59e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X3 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.5425e+11p ps=3.69e+06u w=650000u l=150000u
X4 a_470_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.75e+11p ps=2.55e+06u w=1e+06u l=150000u
X6 a_384_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X7 a_384_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VPWR Y VNB VPB
X0 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=8.3e+11p ps=7.66e+06u w=1e+06u l=150000u
X1 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=1.2415e+12p ps=1.032e+07u w=650000u l=150000u
X2 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X3 a_475_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=8.3e+11p pd=7.66e+06u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X5 VPWR A1 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_475_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y A2 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_2 A VGND VPWR Y VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=2.205e+11p ps=2.73e+06u w=420000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VPWR X VNB VPB
X0 a_429_297# A2 a_345_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=4.3e+11p pd=2.86e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 VGND A2 a_345_47# VNB sky130_fd_pr__nfet_01v8 ad=8.45e+11p pd=6.5e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=150000u
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=1.2e+12p pd=8.4e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X4 a_345_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_345_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_629_297# B2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.8e+11p pd=2.76e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X7 VPWR B1 a_629_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_79_21# B2 a_345_47# VNB sky130_fd_pr__nfet_01v8 ad=2.47e+11p pd=2.06e+06u as=0p ps=0u w=650000u l=150000u
X9 a_345_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_79_21# A3 a_429_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_345_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_8 A VGND VPWR Y VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=4.704e+11p pd=5.6e+06u as=5.754e+11p ps=6.94e+06u w=420000u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=1.875e+12p pd=1.775e+07u as=1.62e+12p ps=1.524e+07u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VPWR X VNB VPB
X0 a_27_47# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1e+12p pd=6e+06u as=9.35e+11p ps=7.87e+06u w=1e+06u l=150000u
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=6.041e+11p pd=5.77e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X2 VPWR C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A1 a_373_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X4 a_182_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=3.4735e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X6 a_182_47# B1 a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_373_297# A2 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_110_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X10 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A1 a_182_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VPWR X VNB VPB
X0 VPWR a_80_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=8.45e+11p pd=7.69e+06u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X1 X a_80_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_80_199# X VNB sky130_fd_pr__nfet_01v8 ad=5.655e+11p pd=5.64e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X3 a_386_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X4 X a_80_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_80_199# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=3.25e+11p pd=2.3e+06u as=0p ps=0u w=650000u l=150000u
X6 a_386_297# B1 a_80_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X7 a_458_47# A1 a_80_199# VNB sky130_fd_pr__nfet_01v8 ad=2.47e+11p pd=2.06e+06u as=0p ps=0u w=650000u l=150000u
X8 VPWR A1 a_386_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A2 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VPWR Y VNB VPB
X0 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.12e+12p pd=1.024e+07u as=1.37e+12p ps=1.274e+07u w=1e+06u l=150000u
X1 a_298_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=3.64e+11p pd=3.72e+06u as=5.98e+11p ps=5.74e+06u w=650000u l=150000u
X2 VGND A1 a_497_47# VNB sky130_fd_pr__nfet_01v8 ad=3.64e+11p pd=3.72e+06u as=7.54e+11p ps=7.52e+06u w=650000u l=150000u
X3 a_664_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=9.05e+11p pd=7.81e+06u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A2 a_497_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_298_47# B1 a_497_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_497_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X9 a_497_47# B1 a_298_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y A2 a_664_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_27_47# C1 a_298_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_497_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR A1 a_664_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_664_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
R0 HI VPWR sky130_fd_pr__res_generic_po w=480000u l=45000u
R1 VGND LO sky130_fd_pr__res_generic_po w=480000u l=45000u
.ends

.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VPWR Y VNB VPB
X0 a_113_297# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=1.94e+12p ps=1.388e+07u w=1e+06u l=150000u
X1 a_113_47# A2_N a_113_297# VNB sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 VPWR B1 a_730_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X3 VPWR A2_N a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_730_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X5 a_471_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=7.1825e+11p pd=7.41e+06u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u
X6 a_471_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y B2 a_730_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_113_297# A2_N a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_113_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A1_N a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND B2 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR a_113_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_113_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y a_113_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_730_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y a_113_297# a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X17 a_471_47# a_113_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR A1_N a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND B1 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2_2 A B VGND VPWR X VNB VPB
X0 X a_61_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=8.307e+11p ps=6.94e+06u w=1e+06u l=150000u
X1 VPWR a_61_75# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR B a_61_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3 VGND B a_147_75# VNB sky130_fd_pr__nfet_01v8 ad=4.706e+11p pd=4.14e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4 X a_61_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=2.535e+11p pd=2.08e+06u as=0p ps=0u w=650000u l=150000u
X5 VGND a_61_75# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_61_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_147_75# A a_61_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VPWR X VNB VPB
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=6.246e+11p ps=6.63e+06u w=420000u l=150000u
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=6.015e+11p pd=5.29e+06u as=0p ps=0u w=420000u l=150000u
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X7 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VPWR Y VNB VPB
X0 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.33e+12p pd=1.266e+07u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X1 a_467_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=5.135e+11p pd=5.48e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X2 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_467_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X4 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=7.9e+11p pd=7.58e+06u as=0p ps=0u w=1e+06u l=150000u
X5 Y A1 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_109_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A2 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=5.135e+11p pd=5.48e+06u as=0p ps=0u w=650000u l=150000u
X10 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt digital_pll clockp[0] clockp[1] dco div[0] div[1] div[2] div[3] div[4] enable
+ ext_trim[0] ext_trim[10] ext_trim[11] ext_trim[12] ext_trim[13] ext_trim[14] ext_trim[15]
+ ext_trim[16] ext_trim[17] ext_trim[18] ext_trim[19] ext_trim[1] ext_trim[20] ext_trim[21]
+ ext_trim[22] ext_trim[23] ext_trim[24] ext_trim[25] ext_trim[2] ext_trim[3] ext_trim[4]
+ ext_trim[5] ext_trim[6] ext_trim[7] ext_trim[8] ext_trim[9] osc resetb VPWR VGND
X_363_ _328_/A _363_/D _318_/X VGND VPWR _363_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_294_ _297_/C _302_/C _301_/A VGND VPWR _294_/X VGND VPWR sky130_fd_sc_hd__or3_2
XFILLER_13_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[1\].id.delayint0 ringosc.dstage\[1\].id.delayen1/Z VGND VPWR ringosc.dstage\[1\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
X_346_ _288_/B ext_trim[3] dco VGND VPWR _346_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_277_ _362_/Q _272_/B _363_/Q _267_/B _226_/B VGND VPWR _359_/D VGND VPWR sky130_fd_sc_hd__a311o_2
X_200_ _196_/A _199_/Y _196_/A _199_/Y VGND VPWR _200_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_2
XFILLER_23_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_329_ _292_/B _232_/B _370_/Q VGND VPWR _329_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[11\].id.delayen1 ringosc.dstage\[11\].id.delayen1/A _331_/X VGND
+ VPWR ringosc.dstage\[11\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
Xringosc.dstage\[10\].id.delayenb0 ringosc.dstage\[10\].id.delayenb1/A _332_/X VGND
+ VPWR ringosc.dstage\[10\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[9\].id.delayenb0 ringosc.dstage\[9\].id.delayenb1/A _334_/X VGND
+ VPWR ringosc.dstage\[9\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
XFILLER_16_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_362_ _328_/A _362_/D _319_/X VGND VPWR _362_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_293_ _367_/Q _221_/B _302_/B _370_/Q _232_/B VGND VPWR _293_/X VGND VPWR sky130_fd_sc_hd__o311a_2
X_276_ _276_/A _276_/B VGND VPWR _360_/D VGND VPWR sky130_fd_sc_hd__or2_2
X_345_ _300_/X ext_trim[17] dco VGND VPWR _345_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_328_ _328_/A VGND VPWR clockp[0] VGND VPWR sky130_fd_sc_hd__buf_2
X_259_ _366_/Q _220_/Y _262_/A VGND _370_/VPB _259_/X VGND _370_/VPB sky130_fd_sc_hd__mux2_1
XFILLER_23_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_87 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[10\].id.delayenb1 ringosc.dstage\[10\].id.delayenb1/A _333_/X VGND
+ VPWR ringosc.dstage\[10\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[9\].id.delayenb1 ringosc.dstage\[9\].id.delayenb1/A _335_/X VGND
+ VPWR ringosc.dstage\[9\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
XFILLER_15_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_361_ _328_/A _361_/D _320_/X VGND VPWR _361_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_292_ _301_/A _292_/B VGND VPWR _299_/B VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_12_34 VGND _370_/VPB VGND _370_/VPB sky130_fd_sc_hd__decap_4
X_275_ _267_/A _267_/B _360_/Q _359_/Q _272_/D VGND VPWR _276_/B VGND VPWR sky130_fd_sc_hd__o221a_2
X_344_ _286_/X ext_trim[4] dco VGND _370_/VPB _344_/X VGND _370_/VPB sky130_fd_sc_hd__mux2_1
XFILLER_23_88 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[4\].id.delayen0 ringosc.dstage\[4\].id.delayen0/A _344_/X VGND _370_/VPB
+ ringosc.dstage\[4\].id.delayen0/Z VGND _370_/VPB sky130_fd_sc_hd__einvp_2
X_327_ _327_/A VGND _370_/VPB _327_/X VGND _370_/VPB sky130_fd_sc_hd__buf_1
X_258_ _262_/A _262_/B VGND VPWR _258_/X VGND VPWR sky130_fd_sc_hd__or2_2
X_189_ _371_/Q _226_/B VGND VPWR _371_/D VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_6_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xringosc.dstage\[10\].id.delaybuf0 ringosc.dstage\[9\].id.delayen0/Z VGND VPWR ringosc.dstage\[10\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[9\].id.delaybuf0 ringosc.dstage\[8\].id.delayen0/Z VGND VPWR ringosc.dstage\[9\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[5\].id.delayenb0 ringosc.dstage\[5\].id.delayenb1/A _342_/X VGND
+ VPWR ringosc.ibufp10/A VGND VPWR sky130_fd_sc_hd__einvn_8
XFILLER_22_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_360_ _328_/A _360_/D _321_/X VGND VPWR _360_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_291_ _369_/Q _368_/Q _367_/Q _370_/Q VGND VPWR _291_/X VGND VPWR sky130_fd_sc_hd__a31o_2
X_274_ _272_/D _268_/A _273_/Y _276_/A VGND VPWR _361_/D VGND VPWR sky130_fd_sc_hd__a31o_2
X_343_ _301_/Y ext_trim[18] dco VGND VPWR _343_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xringosc.dstage\[4\].id.delayen1 ringosc.dstage\[4\].id.delayen1/A _345_/X VGND VPWR
+ ringosc.dstage\[4\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
X_188_ _372_/Q _272_/D _371_/Q _226_/B VGND VPWR _372_/D VGND VPWR sky130_fd_sc_hd__a22o_2
X_257_ _236_/A _251_/X _256_/Y _368_/Q _236_/Y VGND VPWR _368_/D VGND VPWR sky130_fd_sc_hd__a32o_2
X_326_ _370_/Q VGND VPWR _326_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_9_58 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_309_ _327_/A VGND VPWR _309_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_10_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[5\].id.delayenb1 ringosc.dstage\[5\].id.delayenb1/A _343_/X VGND
+ VPWR ringosc.dstage\[5\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[10\].id.delaybuf1 ringosc.dstage\[10\].id.delayenb1/A VGND VPWR ringosc.dstage\[10\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[9\].id.delaybuf1 ringosc.dstage\[9\].id.delayenb1/A VGND VPWR ringosc.dstage\[9\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_13_115 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_290_ _369_/Q _368_/Q _297_/C _370_/Q VGND VPWR _290_/X VGND VPWR sky130_fd_sc_hd__a31o_2
X_273_ _267_/A _267_/B _267_/C VGND VPWR _273_/Y VGND VPWR sky130_fd_sc_hd__o21ai_2
X_342_ _283_/X ext_trim[5] dco VGND VPWR _342_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_187_ _372_/Q _226_/B _373_/Q _272_/D VGND VPWR _373_/D VGND VPWR sky130_fd_sc_hd__a22o_2
X_256_ _256_/A _256_/B VGND VPWR _256_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
X_325_ _327_/A VGND VPWR _325_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_239_ _288_/A _239_/B VGND VPWR _239_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
X_308_ _327_/A VGND VPWR _308_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_19_110 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[5\].id.delaybuf0 ringosc.dstage\[4\].id.delayen0/Z VGND VPWR ringosc.dstage\[5\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_272_ _362_/Q _272_/B _363_/Q _272_/D VGND VPWR _276_/A VGND VPWR sky130_fd_sc_hd__and4_2
Xringosc.dstage\[1\].id.delayenb0 ringosc.dstage\[1\].id.delayenb1/A _350_/X VGND
+ _370_/VPB ringosc.dstage\[1\].id.delayen0/Z VGND _370_/VPB sky130_fd_sc_hd__einvn_8
X_341_ _299_/B ext_trim[19] dco VGND VPWR _341_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xringosc.dstage\[8\].id.delayint0 ringosc.dstage\[8\].id.delayen1/Z VGND VPWR ringosc.dstage\[8\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
XFILLER_4_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_186_ _374_/Q _272_/D _359_/Q _226_/B VGND VPWR _374_/D VGND VPWR sky130_fd_sc_hd__a22o_2
X_255_ _297_/A _236_/A _254_/X VGND VPWR _369_/D VGND VPWR sky130_fd_sc_hd__o21ai_2
X_324_ _327_/A VGND VPWR _324_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_9_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_238_ _224_/A _220_/A _224_/B _237_/X VGND _370_/VPB _262_/A VGND _370_/VPB sky130_fd_sc_hd__o22a_2
X_307_ _327_/A VGND VPWR _307_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_169_ _374_/Q VGND VPWR _193_/B VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_19_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[1\].id.delayenb1 ringosc.dstage\[1\].id.delayenb1/A _351_/X VGND
+ VPWR ringosc.dstage\[1\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[5\].id.delaybuf1 ringosc.dstage\[5\].id.delayenb1/A VGND VPWR ringosc.dstage\[5\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_271_ _362_/Q _272_/B _363_/Q _269_/Y _272_/D VGND VPWR _362_/D VGND VPWR sky130_fd_sc_hd__o221a_2
X_340_ _279_/X ext_trim[6] dco VGND VPWR _340_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xringosc.dstage\[1\].id.delayen0 ringosc.dstage\[1\].id.delayen0/A _350_/X VGND _370_/VPB
+ ringosc.dstage\[1\].id.delayen0/Z VGND _370_/VPB sky130_fd_sc_hd__einvp_2
X_254_ _244_/Y _253_/A _244_/A _253_/Y _236_/Y VGND VPWR _254_/X VGND VPWR sky130_fd_sc_hd__a221o_2
X_185_ _375_/Q _272_/D _360_/Q _226_/B VGND VPWR _375_/D VGND VPWR sky130_fd_sc_hd__a22o_2
X_323_ _327_/A VGND VPWR _323_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_237_ _365_/Q _220_/Y _224_/A _220_/A VGND VPWR _237_/X VGND VPWR sky130_fd_sc_hd__a22o_2
X_306_ _327_/A VGND VPWR _306_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_168_ _359_/Q VGND VPWR _267_/B VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_25_115 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_270_ _164_/Y _269_/Y _226_/B VGND VPWR _363_/D VGND VPWR sky130_fd_sc_hd__a21oi_2
Xringosc.dstage\[1\].id.delayen1 ringosc.dstage\[1\].id.delayen1/A _351_/X VGND VPWR
+ ringosc.dstage\[1\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
X_322_ _327_/A VGND VPWR _322_/X VGND VPWR sky130_fd_sc_hd__buf_1
Xringosc.dstage\[1\].id.delaybuf0 ringosc.dstage\[0\].id.delayen0/Z VGND _370_/VPB
+ ringosc.dstage\[1\].id.delayenb1/A VGND _370_/VPB sky130_fd_sc_hd__clkbuf_2
X_184_ _376_/Q _272_/D _361_/Q _226_/B VGND VPWR _376_/D VGND VPWR sky130_fd_sc_hd__a22o_2
X_253_ _253_/A VGND VPWR _253_/Y VGND VPWR sky130_fd_sc_hd__inv_2
Xringosc.dstage\[4\].id.delayint0 ringosc.dstage\[4\].id.delayen1/Z VGND VPWR ringosc.dstage\[4\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
X_305_ _327_/A VGND VPWR _305_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_236_ _236_/A VGND VPWR _236_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_167_ _360_/Q VGND VPWR _267_/A VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_10_83 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_219_ _219_/A _219_/B VGND VPWR _220_/A VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_25_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_28 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[9\].id.delayen0 ringosc.dstage\[9\].id.delayen0/A _334_/X VGND VPWR
+ ringosc.dstage\[9\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XPHY_2 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xringosc.dstage\[1\].id.delaybuf1 ringosc.dstage\[1\].id.delayenb1/A VGND VPWR ringosc.dstage\[1\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_183_ _377_/Q _272_/D _362_/Q _226_/B VGND VPWR _377_/D VGND VPWR sky130_fd_sc_hd__a22o_2
X_252_ _280_/B _220_/A _251_/X VGND VPWR _253_/A VGND VPWR sky130_fd_sc_hd__o21ai_2
X_321_ _327_/A VGND VPWR _321_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_304_ _288_/A _239_/B _302_/B _370_/Q _232_/B VGND VPWR _304_/X VGND VPWR sky130_fd_sc_hd__o311a_2
X_235_ _301_/A _220_/Y _224_/X _234_/X VGND VPWR _236_/A VGND VPWR sky130_fd_sc_hd__o31a_2
X_166_ _361_/Q VGND VPWR _267_/C VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_1_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_218_ _164_/Y _165_/Y div[4] _216_/B _214_/X VGND VPWR _219_/B VGND VPWR sky130_fd_sc_hd__o221ai_2
Xringosc.dstage\[9\].id.delayen1 ringosc.dstage\[9\].id.delayen1/A _335_/X VGND VPWR
+ ringosc.dstage\[9\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XPHY_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_83 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_182_ dco _182_/B VGND VPWR _327_/A VGND VPWR sky130_fd_sc_hd__nor2_2
X_320_ _327_/A VGND VPWR _320_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_251_ _256_/A _256_/B VGND VPWR _251_/X VGND VPWR sky130_fd_sc_hd__or2_2
X_234_ _219_/B _225_/Y _220_/A _233_/X _226_/X VGND VPWR _234_/X VGND VPWR sky130_fd_sc_hd__o221a_2
X_303_ _297_/A _368_/Q _367_/Q _302_/X VGND VPWR _303_/X VGND VPWR sky130_fd_sc_hd__o31a_2
X_165_ _378_/Q VGND VPWR _165_/Y VGND VPWR sky130_fd_sc_hd__inv_2
Xringosc.iss.reseten0 ringosc.iss.const1/HI _182_/B VGND VPWR ringosc.ibufp00/A VGND
+ VPWR sky130_fd_sc_hd__einvp_1
Xringosc.dstage\[0\].id.delayint0 ringosc.dstage\[0\].id.delayen1/Z VGND VPWR ringosc.dstage\[0\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
X_217_ _201_/Y _203_/Y _205_/Y _211_/Y _216_/Y VGND VPWR _219_/A VGND VPWR sky130_fd_sc_hd__o221a_2
XFILLER_19_83 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[8\].id.delayenb0 ringosc.dstage\[8\].id.delayenb1/A _336_/X VGND
+ VPWR ringosc.dstage\[8\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
XFILLER_23_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_250_ _301_/A _236_/A _249_/X VGND VPWR _370_/D VGND VPWR sky130_fd_sc_hd__o21ai_2
X_181_ enable resetb VGND VPWR _182_/B VGND VPWR sky130_fd_sc_hd__nand2_2
X_302_ _370_/Q _302_/B _302_/C VGND VPWR _302_/X VGND VPWR sky130_fd_sc_hd__and3_2
X_233_ _365_/Q _364_/Q _233_/C VGND VPWR _233_/X VGND VPWR sky130_fd_sc_hd__or3_2
X_164_ _363_/Q VGND VPWR _164_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_216_ div[4] _216_/B VGND VPWR _216_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_18_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xringosc.iss.delayint0 ringosc.iss.delayen1/Z VGND VPWR ringosc.iss.delayen0/A VGND
+ VPWR sky130_fd_sc_hd__clkinv_1
XFILLER_7_54 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_5 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_133 VGND _370_/VPB VGND _370_/VPB sky130_fd_sc_hd__decap_3
Xringosc.dstage\[8\].id.delayenb1 ringosc.dstage\[8\].id.delayenb1/A _337_/X VGND
+ VPWR ringosc.dstage\[8\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
X_180_ _378_/Q _272_/D _363_/Q _226_/B VGND VPWR _378_/D VGND VPWR sky130_fd_sc_hd__a22o_2
X_378_ _328_/A _378_/D _327_/X VGND VPWR _378_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_301_ _301_/A _301_/B VGND VPWR _301_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
X_232_ _370_/Q _232_/B VGND VPWR _233_/C VGND VPWR sky130_fd_sc_hd__or2_2
X_215_ _214_/A _214_/B _214_/X VGND VPWR _216_/B VGND VPWR sky130_fd_sc_hd__a21bo_2
Xringosc.dstage\[6\].id.delayen0 ringosc.dstage\[6\].id.delayen0/A _340_/X VGND VPWR
+ ringosc.dstage\[6\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XPHY_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_377_ _328_/A _377_/D _327_/A VGND VPWR _377_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_1_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[8\].id.delaybuf0 ringosc.dstage\[7\].id.delayen0/Z VGND VPWR ringosc.dstage\[8\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[4\].id.delayenb0 ringosc.dstage\[4\].id.delayenb1/A _344_/X VGND
+ VPWR ringosc.dstage\[4\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
X_300_ _221_/A _366_/Q _301_/A _302_/C _296_/X VGND VPWR _300_/X VGND VPWR sky130_fd_sc_hd__o41a_2
X_231_ _297_/C _302_/B VGND VPWR _232_/B VGND VPWR sky130_fd_sc_hd__or2_2
Xringosc.dstage\[10\].id.delayen0 ringosc.dstage\[10\].id.delayen0/A _332_/X VGND
+ VPWR ringosc.dstage\[10\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
X_214_ _214_/A _214_/B VGND VPWR _214_/X VGND VPWR sky130_fd_sc_hd__or2_2
Xringosc.dstage\[6\].id.delayen1 ringosc.dstage\[6\].id.delayen1/A _341_/X VGND VPWR
+ ringosc.dstage\[6\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XPHY_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_376_ _328_/A _376_/D _305_/X VGND VPWR _376_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[4\].id.delayenb1 ringosc.dstage\[4\].id.delayenb1/A _345_/X VGND
+ _370_/VPB ringosc.dstage\[4\].id.delayen1/Z VGND _370_/VPB sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[8\].id.delaybuf1 ringosc.dstage\[8\].id.delayenb1/A VGND VPWR ringosc.dstage\[8\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_230_ _302_/B VGND VPWR _301_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_359_ _328_/A _359_/D _322_/X VGND VPWR _359_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[10\].id.delayen1 ringosc.dstage\[10\].id.delayen1/A _333_/X VGND
+ VPWR ringosc.dstage\[10\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
X_213_ _362_/Q _377_/Q _190_/Y _376_/Q VGND VPWR _214_/B VGND VPWR sky130_fd_sc_hd__o2bb2a_2
XFILLER_21_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_111 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_8 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_110 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_375_ _328_/A _375_/D _306_/X VGND VPWR _375_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_358_ _328_/A _358_/D _323_/X VGND VPWR _358_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_289_ _297_/A _368_/Q _370_/Q _284_/X VGND VPWR _289_/X VGND VPWR sky130_fd_sc_hd__o31a_2
Xringosc.dstage\[4\].id.delaybuf0 ringosc.dstage\[3\].id.delayen0/Z VGND VPWR ringosc.dstage\[4\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_212_ _363_/Q _378_/Q _164_/Y _165_/Y VGND VPWR _214_/A VGND VPWR sky130_fd_sc_hd__a22o_2
Xringosc.dstage\[0\].id.delayenb0 ringosc.dstage\[0\].id.delayenb1/A _352_/X VGND
+ VPWR ringosc.dstage\[0\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[7\].id.delayint0 ringosc.dstage\[7\].id.delayen1/Z VGND VPWR ringosc.dstage\[7\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
XPHY_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_59 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_68 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_374_ _328_/A _374_/D _307_/X VGND VPWR _374_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_357_ _328_/A _357_/D _324_/X VGND VPWR _358_/D VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_288_ _288_/A _288_/B VGND VPWR _288_/X VGND VPWR sky130_fd_sc_hd__or2_2
Xringosc.dstage\[3\].id.delayen0 ringosc.dstage\[3\].id.delayen0/A _346_/X VGND _370_/VPB
+ ringosc.dstage\[3\].id.delayen0/Z VGND _370_/VPB sky130_fd_sc_hd__einvp_2
X_211_ div[1] _207_/B _210_/X VGND VPWR _211_/Y VGND VPWR sky130_fd_sc_hd__a21oi_2
Xringosc.dstage\[0\].id.delayenb1 ringosc.dstage\[0\].id.delayenb1/A _353_/X VGND
+ VPWR ringosc.dstage\[0\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[4\].id.delaybuf1 ringosc.dstage\[4\].id.delayenb1/A VGND VPWR ringosc.dstage\[4\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xringosc.iss.delayenb0 ringosc.iss.delayenb1/A ringosc.iss.ctrlen0/X VGND VPWR ringosc.ibufp00/A
+ VGND VPWR sky130_fd_sc_hd__einvn_8
XFILLER_16_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_373_ _328_/A _373_/D _308_/X VGND VPWR _373_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_24_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_356_ _328_/A osc _325_/X VGND VPWR _357_/D VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_287_ _297_/A _368_/Q _370_/Q _288_/A _284_/X VGND VPWR _287_/X VGND VPWR sky130_fd_sc_hd__o41a_2
XFILLER_19_68 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xringosc.dstage\[3\].id.delayen1 ringosc.dstage\[3\].id.delayen1/A _347_/X VGND _370_/VPB
+ ringosc.dstage\[3\].id.delayen1/Z VGND _370_/VPB sky130_fd_sc_hd__einvp_2
X_210_ div[1] _207_/B div[0] _209_/Y _207_/Y VGND VPWR _210_/X VGND VPWR sky130_fd_sc_hd__o221a_2
X_339_ _303_/X ext_trim[20] dco VGND VPWR _339_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xringosc.dstage\[0\].id.delaybuf0 ringosc.ibufp00/A VGND VPWR ringosc.dstage\[0\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xringosc.iss.delayenb1 ringosc.iss.delayenb1/A _355_/X VGND VPWR ringosc.iss.delayen1/Z
+ VGND VPWR sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[3\].id.delayint0 ringosc.dstage\[3\].id.delayen1/Z VGND VPWR ringosc.dstage\[3\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
XFILLER_7_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_372_ _328_/A _372_/D _309_/X VGND VPWR _372_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_13_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_286_ _297_/A _368_/Q _370_/Q _367_/Q _284_/X VGND VPWR _286_/X VGND VPWR sky130_fd_sc_hd__o41a_2
X_355_ _304_/X ext_trim[25] dco VGND VPWR _355_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_112 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_269_ _362_/Q _272_/B VGND VPWR _269_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
X_338_ _290_/X ext_trim[7] dco VGND VPWR _338_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xringosc.dstage\[0\].id.delaybuf1 ringosc.dstage\[0\].id.delayenb1/A VGND VPWR ringosc.dstage\[0\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xringosc.iss.delaybuf0 ringosc.iss.delayenb1/A VGND VPWR ringosc.iss.delayen1/A VGND
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_8_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_371_ _328_/A _371_/D _310_/X VGND VPWR _371_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_285_ _297_/A _368_/Q _370_/Q _297_/C _284_/X VGND VPWR _285_/X VGND VPWR sky130_fd_sc_hd__o41a_2
X_354_ _282_/X ext_trim[12] dco VGND VPWR _354_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__diode_2_0 dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_199_ _361_/Q _376_/Q _192_/Y VGND VPWR _199_/Y VGND VPWR sky130_fd_sc_hd__a21oi_2
X_268_ _268_/A VGND VPWR _272_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_337_ _293_/X ext_trim[21] dco VGND VPWR _337_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_116 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_370_ _328_/A _370_/D _311_/X VGND _370_/VPB _370_/Q VGND _370_/VPB sky130_fd_sc_hd__dfrtp_2
XFILLER_24_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_284_ _370_/Q _302_/C _288_/B VGND VPWR _284_/X VGND VPWR sky130_fd_sc_hd__o21a_2
X_353_ _291_/X ext_trim[13] dco VGND VPWR _353_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xringosc.dstage\[0\].id.delayen0 ringosc.dstage\[0\].id.delayen0/A _352_/X VGND VPWR
+ ringosc.dstage\[0\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XFILLER_14_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_198_ _191_/X _376_/Q _191_/X _376_/Q VGND VPWR _202_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_2
X_267_ _267_/A _267_/B _267_/C VGND VPWR _268_/A VGND VPWR sky130_fd_sc_hd__or3_2
Xringosc.dstage\[7\].id.delayenb0 ringosc.dstage\[7\].id.delayenb1/A _338_/X VGND
+ VPWR ringosc.dstage\[7\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
X_336_ _281_/X ext_trim[8] dco VGND VPWR _336_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_25_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_128 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_319_ _327_/A VGND VPWR _319_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_11_131 VGND _370_/VPB VGND _370_/VPB sky130_fd_sc_hd__decap_4
Xringosc.dstage\[0\].id.delayen1 ringosc.dstage\[0\].id.delayen1/A _353_/X VGND VPWR
+ ringosc.dstage\[0\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
X_283_ _370_/Q _302_/C _288_/A _288_/B VGND VPWR _283_/X VGND VPWR sky130_fd_sc_hd__o31a_2
X_352_ _233_/C ext_trim[0] dco VGND VPWR _352_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_197_ _361_/Q _376_/Q _192_/Y _196_/Y VGND VPWR _376_/Q VGND VPWR sky130_fd_sc_hd__o2bb2a_2
X_266_ _364_/Q _236_/A _224_/B _236_/Y VGND VPWR _364_/D VGND VPWR sky130_fd_sc_hd__o22a_2
Xringosc.dstage\[7\].id.delayenb1 ringosc.dstage\[7\].id.delayenb1/A _339_/X VGND
+ VPWR ringosc.dstage\[7\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
X_335_ _296_/X _335_/A1 dco VGND VPWR _335_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_15_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_249_ _246_/Y _248_/A _246_/A _248_/Y _236_/Y VGND _370_/VPB _249_/X VGND _370_/VPB
+ sky130_fd_sc_hd__a221o_2
X_318_ _327_/A VGND _370_/VPB _318_/X VGND _370_/VPB sky130_fd_sc_hd__buf_1
XFILLER_22_83 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[8\].id.delayen0 ringosc.dstage\[8\].id.delayen0/A _336_/X VGND VPWR
+ ringosc.dstage\[8\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XFILLER_5_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_282_ _370_/Q _302_/C _367_/Q _288_/B VGND VPWR _282_/X VGND VPWR sky130_fd_sc_hd__o31a_2
X_351_ _298_/X ext_trim[14] dco VGND _370_/VPB _351_/X VGND _370_/VPB sky130_fd_sc_hd__mux2_1
X_334_ _285_/X ext_trim[9] dco VGND VPWR _334_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_265_ _224_/A _236_/A _236_/Y _264_/X VGND VPWR _365_/D VGND VPWR sky130_fd_sc_hd__o22ai_2
X_196_ _196_/A VGND VPWR _196_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_11_41 VGND _370_/VPB VGND _370_/VPB sky130_fd_sc_hd__decap_4
X_317_ _327_/A VGND VPWR _317_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_248_ _248_/A VGND _370_/VPB _248_/Y VGND _370_/VPB sky130_fd_sc_hd__inv_2
X_179_ _272_/D VGND VPWR _226_/B VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_2_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_52 VGND _370_/VPB VGND _370_/VPB sky130_fd_sc_hd__decap_4
Xringosc.dstage\[7\].id.delaybuf0 ringosc.dstage\[6\].id.delayen0/Z VGND VPWR ringosc.dstage\[7\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[3\].id.delayenb0 ringosc.dstage\[3\].id.delayenb1/A _346_/X VGND
+ VPWR ringosc.dstage\[3\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
XFILLER_20_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[11\].id.delayint0 ringosc.dstage\[11\].id.delayen1/Z VGND VPWR ringosc.dstage\[11\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
Xringosc.dstage\[8\].id.delayen1 ringosc.dstage\[8\].id.delayen1/A _337_/X VGND VPWR
+ ringosc.dstage\[8\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XFILLER_17_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_281_ _297_/C _302_/C _370_/Q _288_/B VGND VPWR _281_/X VGND VPWR sky130_fd_sc_hd__o31a_2
X_350_ _289_/X ext_trim[1] dco VGND VPWR _350_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_264_ _224_/B _237_/X _224_/B _237_/X VGND VPWR _264_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_2
X_195_ _360_/Q _375_/Q _193_/Y _194_/X VGND VPWR _196_/A VGND VPWR sky130_fd_sc_hd__a22o_2
X_333_ _326_/X ext_trim[23] dco VGND VPWR _333_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_84 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_247_ _370_/Q _220_/Y _301_/A _220_/A VGND VPWR _248_/A VGND VPWR sky130_fd_sc_hd__o22a_2
X_316_ _327_/A VGND VPWR _316_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_178_ _358_/D _358_/Q _358_/D _358_/Q VGND VPWR _272_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_2
Xringosc.dstage\[3\].id.delayenb1 ringosc.dstage\[3\].id.delayenb1/A _347_/X VGND
+ _370_/VPB ringosc.dstage\[3\].id.delayen1/Z VGND _370_/VPB sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[7\].id.delaybuf1 ringosc.dstage\[7\].id.delayenb1/A VGND VPWR ringosc.dstage\[7\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_11_101 VGND _370_/VPB VGND _370_/VPB sky130_fd_sc_hd__decap_4
XFILLER_0_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_88 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_280_ _369_/Q _280_/B VGND VPWR _302_/C VGND VPWR sky130_fd_sc_hd__or2_2
X_194_ _360_/Q _375_/Q _360_/Q _375_/Q VGND VPWR _194_/X VGND VPWR sky130_fd_sc_hd__o2bb2a_2
X_263_ _236_/A _258_/X _262_/Y _366_/Q _236_/Y VGND _370_/VPB _366_/D VGND _370_/VPB
+ sky130_fd_sc_hd__a32o_2
X_332_ _288_/X ext_trim[10] dco VGND VPWR _332_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_315_ _327_/A VGND VPWR _315_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_246_ _246_/A VGND VPWR _246_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_177_ div[0] VGND VPWR _177_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_229_ _369_/Q _368_/Q VGND VPWR _302_/B VGND VPWR sky130_fd_sc_hd__or2_2
Xringosc.dstage\[3\].id.delaybuf0 ringosc.dstage\[2\].id.delayen0/Z VGND VPWR ringosc.dstage\[3\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[6\].id.delayint0 ringosc.dstage\[6\].id.delayen1/Z VGND VPWR ringosc.dstage\[6\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
Xringosc.ibufp10 ringosc.ibufp10/A VGND VPWR ringosc.ibufp11/A VGND VPWR sky130_fd_sc_hd__clkinv_2
X_262_ _262_/A _262_/B VGND VPWR _262_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
X_193_ _267_/B _193_/B VGND VPWR _193_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
X_331_ _302_/X ext_trim[24] dco VGND VPWR _331_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_22 VGND _370_/VPB VGND _370_/VPB sky130_fd_sc_hd__decap_3
X_245_ _256_/B _244_/A _256_/A _220_/A _301_/B VGND VPWR _246_/A VGND VPWR sky130_fd_sc_hd__o32a_2
X_314_ _327_/A VGND _370_/VPB _314_/X VGND _370_/VPB sky130_fd_sc_hd__buf_1
X_176_ _364_/Q VGND VPWR _224_/B VGND VPWR sky130_fd_sc_hd__inv_2
Xringosc.dstage\[5\].id.delayen0 ringosc.dstage\[5\].id.delayen0/A _342_/X VGND VPWR
+ ringosc.ibufp10/A VGND VPWR sky130_fd_sc_hd__einvp_2
XFILLER_0_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_54 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_228_ _297_/C VGND VPWR _239_/B VGND VPWR sky130_fd_sc_hd__inv_2
Xringosc.dstage\[3\].id.delaybuf1 ringosc.dstage\[3\].id.delayenb1/A VGND VPWR ringosc.dstage\[3\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_17_54 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_76 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xringosc.ibufp11 ringosc.ibufp11/A VGND VPWR clockp[1] VGND VPWR sky130_fd_sc_hd__clkinv_8
Xringosc.ibufp00 ringosc.ibufp00/A VGND VPWR ringosc.ibufp01/A VGND VPWR sky130_fd_sc_hd__clkinv_2
X_261_ _367_/Q _260_/X _367_/Q _260_/X VGND _370_/VPB _367_/D VGND _370_/VPB sky130_fd_sc_hd__o2bb2a_2
X_192_ _361_/Q _376_/Q VGND VPWR _192_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
X_330_ _287_/X ext_trim[11] dco VGND VPWR _330_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_67 VGND _370_/VPB VGND _370_/VPB sky130_fd_sc_hd__decap_3
X_313_ _327_/A VGND VPWR _313_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_244_ _244_/A VGND VPWR _244_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_175_ _365_/Q VGND VPWR _224_/A VGND VPWR sky130_fd_sc_hd__inv_2
Xringosc.dstage\[5\].id.delayen1 ringosc.dstage\[5\].id.delayen1/A _343_/X VGND VPWR
+ ringosc.dstage\[5\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XFILLER_11_115 VGND _370_/VPB VGND _370_/VPB sky130_fd_sc_hd__decap_4
X_227_ _367_/Q _366_/Q VGND VPWR _297_/C VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_26_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xringosc.dstage\[2\].id.delayint0 ringosc.dstage\[2\].id.delayen1/Z VGND VPWR ringosc.dstage\[2\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
Xringosc.ibufp01 ringosc.ibufp01/A VGND VPWR _328_/A VGND VPWR sky130_fd_sc_hd__clkinv_8
X_260_ _221_/B _220_/A _236_/A _259_/X VGND VPWR _260_/X VGND VPWR sky130_fd_sc_hd__o211a_2
XPHY_22 VGND _370_/VPB VGND _370_/VPB sky130_fd_sc_hd__decap_3
XPHY_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_99 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_191_ _362_/Q _377_/Q _190_/Y VGND VPWR _191_/X VGND VPWR sky130_fd_sc_hd__a21o_2
XFILLER_23_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_243_ _297_/A _220_/Y _369_/Q _220_/A VGND VPWR _244_/A VGND VPWR sky130_fd_sc_hd__o22a_2
X_312_ _327_/A VGND VPWR _312_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_174_ _366_/Q VGND _370_/VPB _221_/B VGND _370_/VPB sky130_fd_sc_hd__inv_2
XFILLER_11_79 VGND _370_/VPB VGND _370_/VPB sky130_fd_sc_hd__decap_6
XFILLER_20_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_226_ _372_/Q _226_/B _373_/Q _371_/Q VGND VPWR _226_/X VGND VPWR sky130_fd_sc_hd__and4_2
Xringosc.dstage\[11\].id.delayenb0 ringosc.dstage\[11\].id.delayenb1/A _330_/X VGND
+ VPWR ringosc.iss.delayenb1/A VGND VPWR sky130_fd_sc_hd__einvn_8
XFILLER_8_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_209_ _209_/A VGND VPWR _209_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_5_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_190_ _362_/Q _377_/Q VGND VPWR _190_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
XPHY_23 VGND _370_/VPB VGND _370_/VPB sky130_fd_sc_hd__decap_3
XPHY_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_242_ _368_/Q _220_/Y _280_/B _220_/A VGND VPWR _256_/B VGND VPWR sky130_fd_sc_hd__a22o_2
X_311_ _327_/A VGND VPWR _311_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_173_ _367_/Q VGND VPWR _221_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_225_ _177_/Y _209_/A _210_/X _205_/A _216_/Y VGND VPWR _225_/Y VGND VPWR sky130_fd_sc_hd__o2111ai_2
Xringosc.dstage\[11\].id.delayenb1 ringosc.dstage\[11\].id.delayenb1/A _331_/X VGND
+ VPWR ringosc.dstage\[11\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
XFILLER_6_110 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_208_ _267_/B _193_/B _193_/Y VGND VPWR _209_/A VGND VPWR sky130_fd_sc_hd__a21oi_2
XFILLER_14_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND _370_/VPB VGND _370_/VPB sky130_fd_sc_hd__decap_3
XPHY_13 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_112 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_310_ _327_/A VGND VPWR _310_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_241_ _239_/Y _262_/B _262_/A _220_/A _239_/B VGND VPWR _256_/A VGND VPWR sky130_fd_sc_hd__o32a_2
Xringosc.iss.const1 VGND VGND VPWR VPWR ringosc.iss.const1/HI ringosc.iss.const1/LO
+ sky130_fd_sc_hd__conb_1
X_172_ _368_/Q VGND VPWR _280_/B VGND VPWR sky130_fd_sc_hd__inv_2
Xringosc.dstage\[2\].id.delayen0 ringosc.dstage\[2\].id.delayen0/A _348_/X VGND VPWR
+ ringosc.dstage\[2\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
X_224_ _224_/A _224_/B _292_/B VGND _370_/VPB _224_/X VGND _370_/VPB sky130_fd_sc_hd__or3_2
XFILLER_12_80 VGND _370_/VPB VGND _370_/VPB sky130_fd_sc_hd__decap_6
XFILLER_17_58 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_207_ div[1] _207_/B VGND VPWR _207_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
Xringosc.dstage\[11\].id.delaybuf0 ringosc.dstage\[10\].id.delayen0/Z VGND VPWR ringosc.dstage\[11\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[6\].id.delayenb0 ringosc.dstage\[6\].id.delayenb1/A _340_/X VGND
+ VPWR ringosc.dstage\[6\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
XFILLER_24_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_25 VGND _370_/VPB VGND _370_/VPB sky130_fd_sc_hd__decap_3
XPHY_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_58 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_240_ _366_/Q _220_/Y _221_/B _220_/A VGND VPWR _262_/B VGND VPWR sky130_fd_sc_hd__a22o_2
X_171_ _369_/Q VGND VPWR _297_/A VGND VPWR sky130_fd_sc_hd__inv_2
Xringosc.dstage\[2\].id.delayen1 ringosc.dstage\[2\].id.delayen1/A _349_/X VGND VPWR
+ ringosc.dstage\[2\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
X_369_ _328_/A _369_/D _312_/X VGND VPWR _369_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_223_ _297_/A _280_/B _223_/C VGND VPWR _292_/B VGND VPWR sky130_fd_sc_hd__or3_2
XFILLER_8_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_206_ _193_/Y _194_/X _193_/Y _194_/X VGND VPWR _207_/B VGND VPWR sky130_fd_sc_hd__o2bb2ai_2
Xringosc.dstage\[6\].id.delayenb1 ringosc.dstage\[6\].id.delayenb1/A _341_/X VGND
+ VPWR ringosc.dstage\[6\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[11\].id.delaybuf1 ringosc.dstage\[11\].id.delayenb1/A VGND VPWR ringosc.dstage\[11\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_5_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_26 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xringosc.iss.delayen0 ringosc.iss.delayen0/A _354_/X VGND VPWR ringosc.ibufp00/A VGND
+ VPWR sky130_fd_sc_hd__einvp_2
X_170_ _370_/Q VGND VPWR _301_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_368_ _328_/A _368_/D _313_/X VGND VPWR _368_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_299_ _329_/X _299_/B VGND VPWR _299_/X VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_9_110 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_222_ _223_/C VGND VPWR _288_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_205_ _205_/A VGND VPWR _205_/Y VGND VPWR sky130_fd_sc_hd__inv_2
Xringosc.dstage\[6\].id.delaybuf0 ringosc.ibufp10/A VGND VPWR ringosc.dstage\[6\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[2\].id.delayenb0 ringosc.dstage\[2\].id.delayenb1/A _348_/X VGND
+ VPWR ringosc.dstage\[2\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[10\].id.delayint0 ringosc.dstage\[10\].id.delayen1/Z VGND VPWR ringosc.dstage\[10\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
Xringosc.dstage\[9\].id.delayint0 ringosc.dstage\[9\].id.delayen1/Z VGND VPWR ringosc.dstage\[9\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
XPHY_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xringosc.iss.delayen1 ringosc.iss.delayen1/A _355_/X VGND VPWR ringosc.iss.delayen1/Z
+ VGND VPWR sky130_fd_sc_hd__einvp_2
X_367_ _328_/A _367_/D _314_/X VGND VPWR _367_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_298_ _301_/A _302_/C _221_/A _297_/X _296_/X VGND VPWR _298_/X VGND VPWR sky130_fd_sc_hd__o311a_2
XFILLER_26_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_221_ _221_/A _221_/B VGND VPWR _223_/C VGND VPWR sky130_fd_sc_hd__or2_2
X_204_ div[2] _200_/X _203_/A _201_/Y VGND VPWR _205_/A VGND VPWR sky130_fd_sc_hd__o211a_2
Xringosc.dstage\[2\].id.delayenb1 ringosc.dstage\[2\].id.delayenb1/A _349_/X VGND
+ VPWR ringosc.dstage\[2\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[6\].id.delaybuf1 ringosc.dstage\[6\].id.delayenb1/A VGND VPWR ringosc.dstage\[6\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_20_83 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_366_ _328_/A _366_/D _315_/X VGND VPWR _366_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_297_ _297_/A _368_/Q _297_/C _301_/A VGND VPWR _297_/X VGND VPWR sky130_fd_sc_hd__or4_2
XFILLER_26_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_220_ _220_/A VGND VPWR _220_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_349_ _295_/X ext_trim[15] dco VGND VPWR _349_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_203_ _203_/A VGND VPWR _203_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_9_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xringosc.iss.ctrlen0 _182_/B _354_/X VGND VPWR ringosc.iss.ctrlen0/X VGND VPWR sky130_fd_sc_hd__or2_2
Xringosc.dstage\[2\].id.delaybuf0 ringosc.dstage\[1\].id.delayen0/Z VGND _370_/VPB
+ ringosc.dstage\[2\].id.delayenb1/A VGND _370_/VPB sky130_fd_sc_hd__clkbuf_2
XPHY_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[5\].id.delayint0 ringosc.dstage\[5\].id.delayen1/Z VGND VPWR ringosc.dstage\[5\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
X_365_ _328_/A _365_/D _316_/X VGND VPWR _365_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_296_ _367_/Q _221_/B _302_/C _301_/A _295_/X VGND VPWR _296_/X VGND VPWR sky130_fd_sc_hd__o41a_2
XFILLER_26_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_96 VGND _370_/VPB VGND _370_/VPB sky130_fd_sc_hd__decap_3
XFILLER_12_52 VGND _370_/VPB VGND _370_/VPB sky130_fd_sc_hd__decap_3
X_279_ _367_/Q _288_/B VGND VPWR _279_/X VGND VPWR sky130_fd_sc_hd__or2_2
X_348_ _284_/X ext_trim[2] dco VGND VPWR _348_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_202_ div[3] _202_/B VGND VPWR _203_/A VGND VPWR sky130_fd_sc_hd__or2_2
Xringosc.dstage\[7\].id.delayen0 ringosc.dstage\[7\].id.delayen0/A _338_/X VGND VPWR
+ ringosc.dstage\[7\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XPHY_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xringosc.dstage\[2\].id.delaybuf1 ringosc.dstage\[2\].id.delayenb1/A VGND _370_/VPB
+ ringosc.dstage\[2\].id.delayen1/A VGND _370_/VPB sky130_fd_sc_hd__clkbuf_1
X_364_ _364_/CLK _364_/D _317_/X VGND VPWR _364_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_295_ _301_/A _302_/B _221_/A _294_/X _293_/X VGND VPWR _295_/X VGND VPWR sky130_fd_sc_hd__o311a_2
XFILLER_13_110 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_278_ _370_/Q _302_/B VGND VPWR _288_/B VGND VPWR sky130_fd_sc_hd__or2_2
X_347_ _299_/X ext_trim[16] dco VGND VPWR _347_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_201_ div[3] _202_/B div[2] _200_/X VGND VPWR _201_/Y VGND VPWR sky130_fd_sc_hd__a22oi_2
XFILLER_9_76 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[11\].id.delayen0 ringosc.dstage\[11\].id.delayen0/A _330_/X VGND
+ VPWR ringosc.iss.delayenb1/A VGND VPWR sky130_fd_sc_hd__einvp_2
Xringosc.dstage\[7\].id.delayen1 ringosc.dstage\[7\].id.delayen1/A _339_/X VGND VPWR
+ ringosc.dstage\[7\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XFILLER_15_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
.ends

